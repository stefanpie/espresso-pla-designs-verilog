module pla__in5 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13;
  assign z00 = (x13 & (((x17 | (~x17 & ~x18)) & ((~x00 & x01 & ((x02 & x03 & x05 & (x07 | (x04 & ~x15))) | (~x02 & x04 & ~x05 & x10 & x11 & x14 & x15 & x16))) | (~x01 & ~x02 & x03 & x04 & ~x05 & ~x09 & x14 & x15 & x16))) | (x04 & ((~x18 & ((~x02 & ~x05 & ((~x01 & x03 & ~x09) | (~x00 & x01 & x10 & x11)) & (~x15 | (x15 & (~x14 | ~x16)))) | (~x00 & x01 & x02 & x03 & x05 & x15))) | (~x00 & x01 & x02 & x03 & x05 & x15 & x17 & (~x14 | ~x16)))) | (~x01 & ~x02 & x03 & x07 & ~x09))) | (~x13 & ~x19 & ~x20 & x21 & x22);
  assign z01 = x13 ? ((~x00 & (x01 ? (x02 ? (x05 & (((x17 ? x15 : ~x18) & (x03 ? x07 : x06)) | (x04 & ((x15 & x16 & (x03 ? (x14 & ~x18) : ~x14)) | (~x17 & ~x18 & ((x03 & (~x14 | ~x15)) | ~x16 | (~x14 & ~x15))))))) : (x04 & ~x05 & x10 & x11 & (x15 ? ((x14 & x16 & (x17 | (~x17 & ~x18))) | (~x18 & (~x14 | ~x16))) : ~x18))) : (x02 & x04 & ~x05 & x10 & (~x16 | (~x14 & (~x15 | (x15 & x16 & (x17 | (~x17 & ~x18))))))))) | (~x01 & ~x02 & ((x04 & ~x05 & ((x15 & ((x16 & (x17 | (~x17 & ~x18)) & ((x03 & ~x09 & x14) | (x00 & ~x03 & ~x14))) | (x03 & ~x09 & ~x18 & (~x14 | ~x16)))) | (x00 & ~x03 & (~x16 | (~x14 & ~x15))) | (x03 & ~x09 & ~x15 & ~x18))) | (x03 & x07 & ~x09) | (x00 & ~x03 & (x06 | x09))))) : (~x21 & x22 & (~x19 ^ x20));
  assign z02 = x13 ? ((~x00 & ((x02 & ((x04 & (((~x16 | (~x14 & ~x15)) & (x01 ? (x05 & (x17 | (~x17 & ~x18))) : (~x05 & x10))) | (x01 & x03 & x05 & ((~x14 & (x17 ? x15 : ~x18)) | (~x15 & (x17 | (~x17 & ~x18))))))) | (x01 & x05 & (x03 ? x07 : x06) & (x17 ? ~x15 : ~x18)))) | (x01 & ~x02 & x04 & ~x05 & x10 & x11 & ~x18 & (~x15 | (x15 & (~x14 | ~x16)))))) | (~x01 & ~x02 & ((x03 & x07 & ~x09) | (x00 & ~x03 & (x06 | x09)) | (x04 & ~x05 & ((x00 & ~x03 & (~x16 | (~x14 & ~x15))) | (x03 & ~x09 & ~x18 & (~x15 | (x15 & (~x14 | ~x16))))))))) : (~x19 & (x20 ? (~x21 & ~x22) : x21));
  assign z03 = (x02 & x13 & ((~x00 & x01 & x05 & (((x17 | (~x17 & ~x18)) & ((x03 & (x07 | (x04 & ~x15))) | (~x03 & x06) | (x04 & ~x14 & ~x15))) | (x04 & ((~x18 & ((x03 & (x14 ? (x15 & x16) : ~x17)) | (~x16 & ~x17))) | (x15 & x16 & ~x03 & ~x14) | (~x15 & ~x16 & x17))))) | (x00 & ~x01 & x03 & x08 & x11))) | (~x13 & x19 & x21 & (x20 ^ x22));
  assign z04 = (x04 & ~x05 & x13 & ((~x02 & ((((~x01 & x03 & ~x09) | (~x00 & x01 & x10 & x11)) & (x15 ? ((~x18 & (~x14 | ~x16)) | (x14 & x16 & x17)) : ~x18)) | (x00 & ~x01 & ~x03 & (~x16 | (~x14 & (~x15 | (x15 & x16 & x17))))))) | (~x00 & ~x01 & x02 & x10 & (~x16 | (~x14 & (~x15 | (x15 & x16 & x17))))))) | (x12 & x18);
  assign z05 = (x12 & x18) | (x04 & x13 & x15 & ((~x05 & ((x16 & (x17 | (~x17 & ~x18)) & ((~x00 & x10 & ((x11 & x14 & x01 & ~x02) | (~x01 & x02 & ~x14))) | (~x01 & ~x02 & ((x03 & ~x09 & x14) | (x00 & ~x03 & ~x14))))) | (~x02 & ((~x18 & ((~x01 & x03 & ~x09) | (~x00 & x01 & x10 & x11)) & (~x14 | ~x16)) | (x00 & ~x01 & ~x03 & ~x16))) | (~x00 & ~x01 & x02 & x10 & ~x16))) | (~x00 & x01 & x02 & x05 & ((x03 & (~x18 | (~x14 & x17))) | (~x16 & (x17 | ~x18)) | (~x03 & ~x14 & x16)))));
  assign z06 = ~x01 & ~x02 & x13 & ((x03 & x07 & ~x09) | (x00 & ~x03 & (x06 | x08 | x09)));
  assign z07 = (x12 & x18) | (x04 & ~x05 & x13 & x15 & ((~x01 & (((~x16 | (~x17 & ~x18 & ~x14 & x16)) & (x00 ? (~x02 & ~x03) : (x02 & x10))) | (~x02 & x03 & ~x09 & ~x18 & (~x14 | ~x16 | (x14 & x16 & ~x17))))) | (~x00 & x01 & ~x02 & x10 & x11 & ~x18 & (~x14 | ~x16 | (x14 & x16 & ~x17)))));
  assign z08 = x13 & ((~x03 & ((x00 & ~x02 & (x08 | (~x01 & (x06 | (x04 & ~x05 & (~x16 | (~x14 & ~x15))))))) | (~x00 & x01 & x02 & ~x17 & ~x18 & x05 & x06))) | (x03 & ((x07 & ((~x01 & ~x02 & ~x09) | (~x00 & x01 & x02 & x05 & ~x17 & ~x18))) | (~x18 & ((x04 & ((~x00 & x01 & x02 & x05 & ~x17 & (~x14 | ~x15)) | (~x01 & ~x02 & ~x05 & ~x09 & (~x15 | (x15 & (~x14 | ~x16)))))) | (~x00 & x01 & x02 & x05 & x23 & (~x14 | ~x15)))))) | (~x00 & ((x01 & ~x02 & x04 & ~x05 & x10 & x11 & ~x18 & (~x15 | (x15 & (~x14 | ~x16)))) | (x02 & (~x16 | (~x14 & ~x15)) & ((x01 & x05 & ~x18 & (x23 | (x04 & ~x17))) | (~x05 & x10 & ~x01 & x04))))));
  assign z09 = x13 & ((x04 & ((x15 & ((x16 & ((~x05 & (x17 | (~x17 & ~x18)) & ((~x00 & x10 & ((x11 & x14 & x01 & ~x02) | (~x01 & x02 & ~x14))) | (~x01 & ~x02 & ((x03 & ~x09 & x14) | (x00 & ~x03 & ~x14))))) | (~x00 & x01 & x02 & x05 & (x03 ? (x14 & ~x18) : ~x14)))) | (~x00 & x01 & x02 & ~x14 & x17 & x03 & x05))) | (~x00 & x01 & x02 & x05 & x17 & (~x16 | (~x15 & (x03 | ~x14)))))) | (~x00 & x01 & x02 & x05 & (x03 ? ((x07 & x17) | (x14 & x15 & x16 & ~x18 & x23)) : ((x06 & x17) | (x16 & ~x18 & x23 & ~x14 & x15)))));
  assign z10 = ~x00 & x04 & ~x05 & x10 & x13 & ((x15 & ((x16 & (x17 | (~x17 & ~x18)) & ((x11 & x14 & x01 & ~x02) | (~x01 & x02 & ~x14))) | (x01 & ~x02 & x11 & ~x18 & (~x14 | ~x16)))) | (~x01 & x02 & (~x16 | (~x14 & ~x15))) | (x01 & ~x02 & x11 & ~x15 & ~x18));
  assign z11 = x13 & x09 & ~x03 & ~x02 & x00 & ~x01;
  assign z12 = x00 & x08 & x13 & (x02 ? ~x01 : ~x03);
  assign z13 = ~x18 & ~x17 & ~x05 & x15;
endmodule