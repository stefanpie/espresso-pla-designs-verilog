module pla__in7 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25,
    z0, z1, z2, z3, z4, z5, z6, z7, z8, z9  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25;
  output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
  assign z0 = x16 | (~x09 & ~x10 & ~x11 & ~x12 & (x13 | (x14 & x15)));
  assign z1 = ((~x21 | x25) & ((x19 & ((~x09 & (x02 | (~x10 & ~x11 & ~x12))) | x00 | (~x01 & x09))) | (~x19 & (~x00 | ~x03 | ~x08)) | ~x15 | x18)) | (((~x18 & x19) | (~x00 & ~x21)) & ((~x09 & (x02 | (~x10 & ~x11 & ~x12))) | x24 | (~x01 & x09))) | (~x18 & (((~x00 | ~x03 | ~x08) & (~x19 | x24)) | ~x15 | x22 | (x00 & x19))) | (~x21 & ((x00 & (~x03 | ~x08)) | (x24 & (~x08 | x19 | (~x03 & ~x25))))) | (x22 & x25);
  assign z2 = (~x00 & ~x09 & ~x18 & x19 & ~x22 & ~x24 & ((~x11 & ((~x02 & x15 & (x10 | (~x10 & x12))) | (~x10 & ~x12 & ~x15 & (x04 | x05 | x06 | x07)))) | (~x02 & x11 & x15))) | (x18 & ~x25);
  assign z3 = x18 ? ~x25 : (~x22 & (x00 ? (x03 & ((~x15 & x19) | (x08 & x15 & ~x19))) : (x19 & ~x24 & ((~x09 & ~x10 & ((~x02 & x15 & (x11 | (~x11 & x12))) | (~x11 & ~x12 & ~x15 & (x06 | x07)))) | (x01 & x09 & x15) | (x02 & ~x15)))));
  assign z4 = (~x18 & ~x22 & (x00 ? (x03 & ((~x15 & x19) | (x08 & x15 & ~x19))) : (x19 & ~x24 & ((x01 & x09 & x15) | (x02 & ~x15) | (~x09 & ~x11 & ((~x02 & x15 & (x10 | (~x10 & x12))) | (~x10 & ~x12 & ~x15 & (x05 | x07)))))))) | (x17 & x18 & ~x25);
  assign z5 = (~x18 & ((~x20 & ~x22 & (x00 ? (x03 & ((x08 & x15 & ~x19) | (~x15 & x19 & ~x23))) : (x19 & ~x24 & ((~x09 & ((~x02 & x15 & (x10 | x11 | x12)) | (~x10 & ~x11 & ~x12 & ~x15 & ~x23 & (x04 | x05 | x06 | x07)))) | (x01 & x09 & x15) | (x02 & ~x15 & ~x23))))) | (x23 & ((~x19 & (~x00 | ~x03 | ~x08)) | ~x15 | x22)))) | (x18 & (x25 ? x23 : ~x20)) | (x23 & (x19 | x20));
  assign z6 = ~x18 & ~x20 & ~x22 & (x00 ? (x03 & ((x08 & x15 & ~x19) | (~x15 & x19 & ~x23))) : (x19 & ~x24 & ((~x09 & ((~x02 & x15 & (x10 | x11 | x12)) | (~x10 & ~x11 & ~x12 & ~x15 & ~x23 & (x04 | x05 | x06 | x07)))) | (x01 & x09 & x15) | (x02 & ~x15 & ~x23))));
  assign z7 = ~x25 & x18 & ~x20;
  assign z8 = x23 & ((~x18 & ((~x19 & (~x00 | ~x03 | ~x08)) | ~x15 | x22 | (x19 & ((~x09 & (x02 | (~x10 & ~x11 & ~x12))) | x00 | x24 | (~x01 & x09))))) | x20 | (x18 & x25));
  assign z9 = x12 & ~x11 & ~x09 & ~x10;
endmodule