module pla__ibm ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    x42, x43, x44, x45, x46, x47,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    x41, x42, x43, x44, x45, x46, x47;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16;
  assign z00 = (x07 & ((x06 & ((~x08 & ((x04 & (((x03 | x09) & ((x00 & x01 & x02 & ~x05) | (~x02 & x05 & x12 & x13))) | (x02 & x05 & ((x09 & x11) | (~x03 & ~x09 & x12))))) | (x15 & (~x04 | (~x05 & (~x02 | (~x03 & ~x09))))))) | (x02 & x03 & x04 & x05 & ~x10 & x11) | (~x04 & ~x05 & x08 & ~x16))) | (~x04 & x05 & ~x08 & x15))) | (x14 & ((x00 & x01 & x02 & (x03 | x09)) | (x15 & (~x02 | (~x03 & ~x09))))) | (~x04 & ~x05 & ~x06 & ~x07 & x15);
  assign z01 = ((x03 | x09) & (((x14 | (~x04 & ~x05 & x06 & x07 & x08 & ~x16)) & (x02 ? x11 : (x12 & x13))) | (x02 & x04 & ~x05 & x06 & x07 & ~x08 & x11))) | (~x03 & ~x09 & ((x02 & x12 & (x14 | (~x04 & ~x05 & x06 & x07 & x08 & ~x16))) | (~x05 & x06 & x07 & ~x08 & x17))) | (x07 & x17 & ((~x04 & (x05 ? ~x08 : x06)) | (~x02 & ~x05 & x06 & ~x08)));
  assign z02 = ((x14 | (x04 & x06 & x07 & ~x08)) & ((x18 & (~x02 | (~x03 & ~x09) | (~x16 & (~x00 | ~x01)))) | (x16 & x19))) | (~x04 & x18 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z03 = ((x14 | (x04 & x06 & x07 & ~x08)) & ((x20 & (~x02 | (~x03 & ~x09) | (~x00 & ~x16))) | (x16 & x21))) | (x20 & ((~x01 & ((x04 & x06 & x07 & ~x08 & x16) | (x14 & ~x16))) | (~x04 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)))));
  assign z04 = (x22 & ((~x00 & ((x04 & x06 & x07 & ~x08 & x16) | (x14 & ~x16))) | (~x04 & (x05 ? (x07 & ~x08) : (~x06 ^ x07))) | ((x14 | (x04 & x06 & x07 & ~x08)) & (~x02 | (~x03 & ~x09) | (~x01 & ~x16))))) | (x16 & x23 & (x14 | (x04 & x06 & x07 & ~x08)));
  assign z05 = ((x14 | (x04 & x06 & x07 & ~x08)) & ((x24 & (~x02 | (~x03 & ~x09) | (~x16 & (~x00 | ~x01)))) | (x16 & x25))) | (~x04 & x24 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z06 = (x26 & ((~x16 & ((~x00 & (x14 | (x07 & ~x08 & x04 & x05))) | (~x01 & (x14 | (x04 & x06 & x07 & ~x08))))) | ((~x02 | (~x03 & ~x09)) & (x14 | (x04 & x06 & x07 & ~x08))) | (~x04 & ~x05 & (x07 ? (x06 | ~x08) : ~x06)))) | (x16 & x27 & (x14 | (x04 & x06 & x07 & ~x08)));
  assign z07 = ((x14 | (x04 & x06 & x07 & ~x08)) & ((x28 & (~x02 | (~x03 & ~x09) | (~x16 & (~x00 | ~x01)))) | (x16 & x29))) | (~x04 & x28 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z08 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x31 : x30)) | (~x04 & x07 & x30 & (x05 ? ~x08 : ~x06));
  assign z09 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x33 : x32)) | (~x04 & x32 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z10 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x35 : x34)) | (~x04 & x34 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z11 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x37 : x36)) | (~x04 & x36 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z12 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x39 : x38)) | (~x04 & x38 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z13 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x41 : x40)) | (~x04 & x40 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z14 = (x07 & ((x06 & (x04 ? (~x08 & (x16 ? x43 : x42)) : (~x05 & x42))) | (~x04 & x05 & ~x08 & x42))) | (x14 & (x16 ? x43 : x11)) | (~x04 & ~x05 & ~x06 & ~x07 & x42);
  assign z15 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x45 : x44)) | (~x04 & x44 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
  assign z16 = ((x14 | (x04 & x06 & x07 & ~x08)) & (x16 ? x47 : x46)) | (~x04 & x46 & (x05 ? (x07 & ~x08) : (~x06 ^ x07)));
endmodule