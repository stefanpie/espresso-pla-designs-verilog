module pla__exep ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62;
  assign z00 = (~x01 & (x00 ? (x02 ? ((~x12 & ((x03 & x04 & x13 & x15) | (~x03 & ~x04 & ~x13 & x14 & ~x15 & ~x16))) | (x12 & ((x03 & x04 & (~x14 | ~x15)) | (~x03 & ~x04 & ~x13 & ~x15))) | (~x03 & ~x04 & ~x16 & (x13 ? (~x14 | (x14 & ~x15)) : (x14 & x15)))) : ((x04 & (x03 ? (~x07 & ((~x06 & (~x05 | (x05 & ~x14 & ~x16))) | (~x05 & x06 & x08 & x09 & x10 & ~x16 & (x11 ? (~x12 | (x12 & (x13 ^ x14))) : x12)))) : (~x11 & (x12 | (~x12 & (~x14 | x15 | (x14 & ~x15))))))) | (~x03 & ~x04 & (x11 ? ~x12 : ((x12 & (x13 ? ~x15 : (x14 & ~x16))) | (~x13 & (~x14 | (~x12 & x14))) | (x13 & x15 & ~x16 & (x14 | (~x14 & (x07 | (x06 & ~x07))))) | (~x14 & ~x15)))))) : ((~x13 & ((x02 & ~x03 & x04) | (~x02 & x03 & ~x04 & ~x12))) | (x02 & ~x03 & (~x04 | (x04 & (x12 | (x14 & x15 & ~x12 & x13))))) | (~x02 & x03 & ~x04 & ((x12 & (~x14 ^ ~x15)) | (x13 & ((x14 & ~x15) | (~x12 & ~x14 & x15)))))))) | (x01 & ((x03 & (x00 ? (~x02 & (x04 | (~x04 & ((~x05 & ~x06 & ~x07) | (x14 & ~x15) | (~x08 & ~x09 & ~x10))))) : (x02 ? (~x14 | ~x15) : ~x04))) | (~x02 & ~x03 & (x00 ? (~x04 | (x04 & (~x13 | (x13 & x14 & ~x15)))) : x04)))) | (~x00 & x02 & ~x03 & x04 & (~x14 | ~x15));
  assign z01 = x20 & x22 & x23 & x24 & x25 & x27 & ((~x04 & (x00 ? (~x01 & ~x02 & x03 & x12 & (~x13 | x14 | x15 | (x13 & ~x14 & ~x15))) : (~x03 & (x01 | (~x01 & ~x02))))) | (x00 & x02 & ~x03 & (x01 | (~x01 & x04))));
  assign z02 = ~x01 & x03 & x20 & x22 & x26 & x27 & ((x04 & ((~x00 & ~x02) | (~x13 & x14 & x15 & x00 & x02 & x12))) | ((x13 | ~x14) & ((~x00 & x02 & x12) | (~x04 & ~x12 & x00 & ~x02))));
  assign z03 = x03 & x20 & x22 & x25 & x26 & x29 & ((~x00 & (x01 ? (~x02 & x04) : (x02 & ~x12 & (x13 | ~x14)))) | (~x02 & ~x04 & x00 & ~x01 & x14 & ~x15 & ~x12 & ~x13));
  assign z04 = x00 & ~x01 & x02 & x03 & x04 & x20 & x22 & x24 & x25 & x26 & x29 & ((~x12 & (~x13 | (x14 & ~x15))) | (x14 & x15 & x12 & x13));
  assign z05 = x00 & ~x01 & ~x03 & ~x04 & ~x06 & x07 & x12 & x13 & ~x14 & x15 & ~x16 & x19 & x22 & x26 & x28 & x29 & (x02 | (~x02 & ~x11));
  assign z06 = x00 & ~x01 & ~x14 & ~x15 & x20 & x21 & x22 & x24 & x25 & x26 & x29 & ((x02 & x03 & x04 & ~x12 & x13) | (~x02 & ~x03 & ~x04 & x11 & x12 & ~x13));
  assign z07 = x00 & x01 & ~x02 & ~x03 & x04 & x13 & x20 & x21 & x23 & x24 & x26 & x28 & x29 & (x14 | x15);
  assign z08 = x00 & ~x01 & ~x03 & ~x04 & x06 & x07 & x12 & x13 & ~x14 & x15 & ~x16 & x21 & x22 & x23 & x24 & x26 & x28 & x29 & (x02 | (~x02 & ~x11));
  assign z09 = x00 & ~x01 & ~x03 & ~x04 & ~x06 & ~x07 & x12 & x13 & ~x14 & x15 & ~x16 & x21 & x22 & x23 & x24 & x26 & x29 & (x02 | (~x02 & ~x11));
  assign z10 = x00 & ~x01 & ~x03 & ~x04 & x06 & ~x07 & x12 & x13 & ~x14 & x15 & ~x16 & x22 & x23 & x26 & x29 & (x02 | (~x02 & ~x11));
  assign z11 = x28 & x23 & x22 & x21 & x20 & x19 & x07 & x06 & x05 & x04 & x03 & ~x02 & x00 & ~x01;
  assign z12 = x29 & x27 & x25 & x24 & x22 & x21 & x20 & x19 & ~x15 & ~x14 & x12 & ~x04 & x03 & ~x02 & x00 & x01;
  assign z13 = x29 & x28 & x27 & x24 & x22 & x21 & x20 & x19 & x15 & ~x14 & x12 & ~x04 & x03 & ~x02 & x00 & x01;
  assign z14 = x29 & x28 & x26 & x23 & x21 & x20 & x19 & x15 & x14 & ~x13 & x12 & ~x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z15 = x29 & x28 & x27 & x23 & x21 & x20 & x19 & x15 & x14 & x13 & x12 & ~x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z16 = x29 & x27 & x26 & x21 & x20 & x19 & ~x16 & x09 & ~x08 & ~x07 & x06 & ~x05 & x04 & x03 & ~x02 & x00 & ~x01;
  assign z17 = x29 & x27 & x21 & x20 & x19 & ~x16 & ~x09 & ~x08 & ~x07 & x06 & ~x05 & x04 & x03 & ~x02 & x00 & ~x01;
  assign z18 = x29 & x28 & x25 & x24 & x23 & x22 & x20 & x19 & x15 & ~x14 & x13 & ~x12 & x04 & x03 & x02 & x00 & ~x01;
  assign z19 = x29 & x28 & x26 & x22 & x20 & x19 & ~x15 & ~x14 & ~x13 & x12 & ~x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z20 = x29 & x28 & x22 & x20 & x19 & ~x15 & ~x14 & x13 & x12 & ~x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z21 = x29 & x28 & x27 & x26 & x25 & x24 & x23 & x20 & x19 & ~x16 & x15 & ~x14 & ~x13 & ~x12 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z22 = x27 & x25 & x23 & x20 & x19 & ~x16 & x15 & x14 & ~x13 & ~x12 & x07 & ~x06 & x05 & ~x04 & x03 & ~x02 & x00 & ~x01;
  assign z23 = x27 & x26 & x23 & x20 & x19 & x15 & x14 & x13 & ~x12 & x04 & x03 & x02 & x00 & ~x01;
  assign z24 = x27 & x25 & x24 & x20 & x19 & ~x16 & x15 & x14 & ~x13 & ~x12 & x07 & x06 & ~x04 & x03 & ~x02 & x00 & ~x01;
  assign z25 = x27 & x25 & x20 & x19 & ~x16 & x15 & x14 & ~x13 & ~x12 & ~x07 & ~x04 & x03 & ~x02 & x00 & ~x01;
  assign z26 = x26 & x22 & x21 & x19 & ~x16 & x15 & ~x14 & x13 & ~x12 & x07 & ~x06 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z27 = x28 & x25 & x24 & x23 & x21 & x19 & x15 & ~x14 & ~x12 & ~x04 & x03 & ~x02 & x00 & x01;
  assign z28 = x29 & x24 & x23 & x21 & x19 & x14 & x12 & ~x04 & x03 & ~x02 & x00 & x01;
  assign z29 = x26 & x23 & x21 & x19 & ~x16 & x15 & ~x14 & x13 & ~x12 & ~x07 & ~x06 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z30 = x28 & x27 & x25 & x24 & x21 & x19 & ~x15 & ~x14 & ~x12 & ~x04 & x03 & ~x02 & x00 & x01;
  assign z31 = x29 & x28 & x27 & x26 & x24 & x21 & x19 & x15 & x14 & ~x12 & ~x04 & x03 & ~x02 & x00 & x01;
  assign z32 = x29 & x26 & x21 & x19 & ~x16 & x15 & ~x14 & x13 & ~x12 & x07 & x06 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z33 = x26 & x22 & x19 & ~x16 & x15 & ~x14 & x13 & ~x12 & ~x07 & x06 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z34 = x28 & x27 & x26 & x25 & x24 & x23 & x19 & x17 & x15 & x14 & x13 & ~x12 & x04 & ~x03 & x02 & ~x00 & x01;
  assign z35 = x28 & x27 & x26 & x24 & x23 & x19 & x17 & x15 & x14 & ~x13 & ~x12 & x04 & ~x03 & x02 & ~x00 & x01;
  assign z36 = x28 & x27 & x26 & x25 & x24 & x19 & ~x17 & x15 & x14 & x13 & ~x12 & x04 & ~x03 & x02 & ~x00 & x01;
  assign z37 = x28 & x27 & x26 & x24 & x19 & ~x17 & x15 & x14 & ~x13 & ~x12 & x04 & ~x03 & x02 & ~x00 & x01;
  assign z38 = x28 & x27 & x26 & x25 & x19 & x15 & x14 & ~x13 & x12 & x04 & ~x03 & x02 & ~x00 & x01;
  assign z39 = x28 & x27 & x26 & x19 & x15 & x14 & x13 & x12 & x04 & ~x03 & x02 & ~x00 & x01;
  assign z40 = x29 & x28 & x27 & x26 & x22 & x21 & x20 & ~x15 & ~x14 & x13 & ~x12 & ~x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z41 = x29 & x28 & x27 & x26 & x23 & x21 & x20 & x15 & x14 & x13 & ~x12 & ~x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z42 = x28 & x27 & x26 & x25 & x24 & x23 & x22 & x20 & ~x16 & x15 & x14 & x13 & x12 & x07 & x06 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z43 = x29 & x26 & x25 & x24 & x23 & x22 & x20 & x07 & x06 & ~x05 & x04 & x03 & ~x02 & x00 & ~x01;
  assign z44 = x29 & x27 & x25 & x24 & x23 & x22 & x20 & ~x16 & x15 & x14 & x13 & ~x12 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z45 = x28 & x25 & x24 & x23 & x22 & x20 & ~x16 & ~x15 & ~x14 & ~x13 & ~x12 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z46 = x28 & x26 & x25 & x24 & x20 & ~x16 & x14 & x13 & x12 & x11 & x10 & x09 & x08 & ~x07 & x06 & ~x05 & x04 & x03 & ~x02 & x00 & ~x01;
  assign z47 = x29 & x26 & x25 & x20 & x15 & x14 & ~x13 & x03 & x02 & ~x00 & ~x01;
  assign z48 = x28 & x27 & x25 & x20 & ~x16 & x15 & ~x14 & ~x13 & x12 & ~x04 & ~x03 & x02 & x00 & ~x01;
  assign z49 = x28 & x25 & x20 & ~x16 & ~x07 & x06 & x05 & x04 & x03 & ~x02 & x00 & ~x01;
  assign z50 = x26 & x20 & ~x15 & x14 & ~x13 & x03 & x02 & ~x00 & ~x01;
  assign z51 = x27 & x26 & x25 & x24 & x23 & x17 & x15 & x14 & x13 & ~x12 & x03 & x02 & ~x00 & x01;
  assign z52 = x27 & x26 & x24 & x23 & x17 & x15 & x14 & ~x13 & ~x12 & x03 & x02 & ~x00 & x01;
  assign z53 = x27 & x26 & x25 & x23 & x15 & x14 & ~x13 & x12 & x04 & x03 & x02 & ~x00 & x01;
  assign z54 = x27 & x26 & x25 & x24 & ~x17 & x15 & x14 & x13 & ~x12 & x03 & x02 & ~x00 & x01;
  assign z55 = x27 & x26 & x24 & ~x17 & x15 & x14 & ~x13 & ~x12 & x03 & x02 & ~x00 & x01;
  assign z56 = x27 & x26 & x25 & x15 & x14 & ~x13 & x12 & ~x04 & x03 & x02 & ~x00 & x01;
  assign z57 = x27 & x26 & x15 & x14 & x13 & x12 & x03 & x02 & ~x00 & x01;
  assign z58 = x29 & x27 & ~x16 & x15 & ~x14 & x13 & ~x12 & ~x11 & ~x07 & x06 & ~x04 & ~x03 & ~x02 & x00 & ~x01;
  assign z59 = x27 & ~x16 & x15 & ~x14 & x13 & ~x12 & ~x11 & x07 & ~x06 & ~x04 & ~x03 & ~x02 & x00 & ~x01;
  assign z60 = x28 & ~x16 & x15 & ~x14 & x13 & ~x12 & ~x11 & x07 & x06 & ~x04 & ~x03 & ~x02 & x00 & ~x01;
  assign z61 = x29 & ~x16 & x15 & ~x14 & x13 & ~x12 & ~x11 & ~x07 & ~x06 & ~x04 & ~x03 & ~x02 & x00 & ~x01;
  assign z62 = 1'b0;
endmodule