module pla__newcpla1 ( 
    WAIT, CPIPE1s__larrow__0__rarrow__, CPIPE1s__larrow__1__rarrow__,
    CPIPE1s__larrow__2__rarrow__, CPIPE1s__larrow__3__rarrow__,
    CPIPE1s__larrow__4__rarrow__, CPIPE1s__larrow__5__rarrow__,
    CPIPE1s__larrow__7__rarrow__, RESET,
    changeCWP2t, trap, lastPCload, pDATABUSintoLOADL, enableINTS1,
    changeCWP1, PCtoMAL1, pALUtoMAL, pPCIncr, pALUtoPC, DST2step1,
    PCstuffoncall1, SRC2smin1, DST1min1, CPIPE1flush, CPIPE1load1  );
  input  WAIT, CPIPE1s__larrow__0__rarrow__,
    CPIPE1s__larrow__1__rarrow__, CPIPE1s__larrow__2__rarrow__,
    CPIPE1s__larrow__3__rarrow__, CPIPE1s__larrow__4__rarrow__,
    CPIPE1s__larrow__5__rarrow__, CPIPE1s__larrow__7__rarrow__, RESET;
  output changeCWP2t, trap, lastPCload, pDATABUSintoLOADL, enableINTS1,
    changeCWP1, PCtoMAL1, pALUtoMAL, pPCIncr, pALUtoPC, DST2step1,
    PCstuffoncall1, SRC2smin1, DST1min1, CPIPE1flush, CPIPE1load1;
  assign changeCWP2t = CPIPE1s__larrow__7__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~WAIT & CPIPE1s__larrow__0__rarrow__;
  assign trap = CPIPE1s__larrow__7__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__;
  assign lastPCload = ~WAIT & ((CPIPE1s__larrow__7__rarrow__ & ((~CPIPE1s__larrow__3__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__4__rarrow__) | (CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | ~CPIPE1s__larrow__2__rarrow__ | (CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & (CPIPE1s__larrow__1__rarrow__ | (~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__3__rarrow__))))) | CPIPE1s__larrow__5__rarrow__ | (~CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__7__rarrow__));
  assign pDATABUSintoLOADL = ~WAIT & ((CPIPE1s__larrow__0__rarrow__ & (~CPIPE1s__larrow__5__rarrow__ | (~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__))) | (CPIPE1s__larrow__7__rarrow__ & ((CPIPE1s__larrow__1__rarrow__ & ((~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | (~CPIPE1s__larrow__1__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | (~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & (~CPIPE1s__larrow__5__rarrow__ | (CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__5__rarrow__))))) | ~CPIPE1s__larrow__4__rarrow__ | ~CPIPE1s__larrow__7__rarrow__);
  assign enableINTS1 = CPIPE1s__larrow__7__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__;
  assign changeCWP1 = ~CPIPE1s__larrow__7__rarrow__ & ~WAIT & ~CPIPE1s__larrow__5__rarrow__;
  assign PCtoMAL1 = ~WAIT & CPIPE1s__larrow__7__rarrow__ & ((~CPIPE1s__larrow__3__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__4__rarrow__) | (CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | (CPIPE1s__larrow__5__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & (~CPIPE1s__larrow__4__rarrow__ | (~CPIPE1s__larrow__1__rarrow__ & ~CPIPE1s__larrow__2__rarrow__))) | (~CPIPE1s__larrow__4__rarrow__ & (CPIPE1s__larrow__1__rarrow__ ? (CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__3__rarrow__) : (~CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__))))));
  assign pALUtoMAL = ~WAIT & ((CPIPE1s__larrow__0__rarrow__ & ((CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__))) | (CPIPE1s__larrow__7__rarrow__ & ((CPIPE1s__larrow__2__rarrow__ & ((CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | (CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__))) | ~CPIPE1s__larrow__7__rarrow__ | (~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__5__rarrow__));
  assign pPCIncr = ~WAIT & CPIPE1s__larrow__7__rarrow__ & ~RESET & ((CPIPE1s__larrow__5__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & (~CPIPE1s__larrow__4__rarrow__ | (~CPIPE1s__larrow__1__rarrow__ & ~CPIPE1s__larrow__2__rarrow__))) | (~CPIPE1s__larrow__4__rarrow__ & (CPIPE1s__larrow__1__rarrow__ ? (CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__3__rarrow__) : (~CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__))))) | (~CPIPE1s__larrow__3__rarrow__ & ((CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__) | (CPIPE1s__larrow__2__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__4__rarrow__) | (~CPIPE1s__larrow__1__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))))));
  assign pALUtoPC = ~WAIT & ~RESET & (~CPIPE1s__larrow__7__rarrow__ | (CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__));
  assign DST2step1 = ~WAIT & (CPIPE1s__larrow__5__rarrow__ | (CPIPE1s__larrow__7__rarrow__ & ((~CPIPE1s__larrow__3__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__4__rarrow__) | (CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | ~CPIPE1s__larrow__2__rarrow__ | (CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & (CPIPE1s__larrow__1__rarrow__ | (~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__3__rarrow__))))));
  assign PCstuffoncall1 = ~CPIPE1s__larrow__7__rarrow__ & ~WAIT & ~CPIPE1s__larrow__5__rarrow__;
  assign SRC2smin1 = ~WAIT & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__7__rarrow__ & ((CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (CPIPE1s__larrow__1__rarrow__ & (CPIPE1s__larrow__5__rarrow__ | (~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__2__rarrow__))));
  assign DST1min1 = ~WAIT & ~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__ & (CPIPE1s__larrow__0__rarrow__ | CPIPE1s__larrow__1__rarrow__ | CPIPE1s__larrow__2__rarrow__);
  assign CPIPE1flush = ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__ & ~RESET & (CPIPE1s__larrow__3__rarrow__ | (CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__2__rarrow__));
  assign CPIPE1load1 = ~WAIT & ~RESET & (~CPIPE1s__larrow__4__rarrow__ | ~CPIPE1s__larrow__5__rarrow__ | ~CPIPE1s__larrow__7__rarrow__);
endmodule