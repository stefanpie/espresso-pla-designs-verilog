module pla__ex5 ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62;
  assign z00 = ~x6 & ~x4 & ~x5;
  assign z01 = ~x7 & ~x5 & ~x6;
  assign z02 = ~x7 & ~x6 & x5 & ~x3 & ~x4;
  assign z03 = ~x7 & ~x6 & x5 & x3 & ~x4;
  assign z04 = ~x7 & x6 & ~x5 & x3 & ~x4;
  assign z05 = ~x7 & x6 & ~x4 & x5;
  assign z06 = ~x6 & ~x5 & ~x4 & x3 & x2 & ~x0 & ~x1;
  assign z07 = x7 & x6 & x5 & ~x4 & ~x3 & ~x2 & ~x0 & x1;
  assign z08 = x7 & x6 & x5 & ~x4 & ~x3 & x2 & x0 & x1;
  assign z09 = x7 & x6 & ~x5 & ~x4 & ~x3 & x2 & ~x0 & ~x1;
  assign z10 = x7 & x6 & x5 & ~x4 & x2 & ~x0 & x1;
  assign z11 = x7 & x6 & x5 & ~x4 & ~x3 & ~x2 & x0 & x1;
  assign z12 = x7 & x6 & x5 & ~x4 & ~x3 & x2 & x0 & ~x1;
  assign z13 = x7 & x6 & x5 & ~x4 & x3 & ~x2 & ~x0 & x1;
  assign z14 = x7 & x6 & x5 & ~x4 & x3 & ~x2 & x0 & ~x1;
  assign z15 = x7 & x6 & x5 & ~x4 & x3 & x2 & ~x0 & x1;
  assign z16 = x7 & x6 & x5 & ~x4 & x3 & ~x2 & x0 & x1;
  assign z17 = ~x5 & x4 & ~x2 & x0 & ~x1;
  assign z18 = ~x5 & x4 & x3 & x2 & ~x0 & ~x1;
  assign z19 = x4 & ~x3 & ~x2 & ~x0 & ~x1;
  assign z20 = ~x6 & ~x5 & ~x4 & ~x3 & ~x2 & x0 & ~x1;
  assign z21 = ~x6 & ~x5 & ~x4 & x3 & ~x2 & x0 & ~x1;
  assign z22 = x7 & x6 & ~x5 & ~x4 & ~x2 & x0 & ~x1;
  assign z23 = x5 & x3 & ~x2 & ~x0 & ~x1;
  assign z24 = ~x7 & x6 & ~x5 & ~x4 & ~x3 & ~x2 & ~x0 & ~x1;
  assign z25 = ~x7 & x6 & ~x5 & ~x4 & ~x3 & ~x2 & ~x0 & x1;
  assign z26 = x7 & x6 & ~x5 & ~x4 & ~x3 & x0 & x2;
  assign z27 = ~x7 & x6 & ~x5 & ~x4 & ~x3 & x2 & ~x0 & x1;
  assign z28 = x7 & x6 & ~x5 & ~x4 & x3 & x2 & x0 & ~x1;
  assign z29 = x7 & ~x6 & ~x5 & ~x4 & ~x3 & ~x2 & ~x0 & ~x1;
  assign z30 = x7 & x6 & ~x5 & ~x4 & ~x3 & x2 & x0 & x1;
  assign z31 = (((x1 & (~x2 | (x0 & x2))) | (~x0 & x2)) & (~x3 | (x3 & (~x4 | (x4 & ~x5))))) | (~x2 & ((~x0 & ((~x1 & ~x4) | (x3 & x4 & x5))) | (x4 & ((x0 & x1 & x3 & x5) | (~x1 & ~x5))) | (x0 & ~x1 & ~x4 & (x6 | (x5 & ~x6))))) | (x2 & ((x0 & ~x1) | (x4 & x5 & x1 & x3)));
  assign z32 = (~x0 & ((~x2 & ((~x1 & (((~x6 | (x6 & x7)) & (x4 ? x5 : ~x3)) | (~x3 & x5 & x6 & ~x7))) | (x3 & x4 & x5 & x6 & ~x7))) | (x3 & (~x4 | (x1 & x4 & (~x5 | (x5 & (~x6 | (x6 & x7))))))) | (x2 & ~x3))) | (x0 & ((x3 & ((~x2 & (x1 | (~x1 & ~x4 & x6))) | (x2 & ((x4 & ((x5 & ~x6) | (x1 & (~x5 | (x5 & x6 & x7))))) | (~x1 & (~x5 | (x5 & x6))))) | (~x1 & ~x4 & x5 & ~x6))) | (x2 & (x4 ? ~x3 : x1)) | (~x1 & ~x3 & ~x4))) | (x1 & ((~x2 & ~x3) | (x5 & x6 & ~x7 & x2 & x3 & x4))) | (x4 & ~x5 & ~x1 & ~x2);
  assign z33 = ~x0 | (x0 & (~x2 | (x2 & (((x1 ? x3 : x4) & (~x5 | (x5 & (~x6 | (x6 & ~x7))))) | (x1 & ((x4 & (~x3 | (x3 & x5 & x6 & x7))) | (~x3 & ~x4 & (~x6 | (x6 & ~x7))))) | (~x1 & ((x5 & x6 & x7) | (~x4 & (~x6 | (x6 & ~x7)))))))));
  assign z34 = (x2 & ((~x0 & ((~x5 & (x4 | (x3 & ~x4))) | (~x3 & (((~x6 | (x6 & x7)) & (x4 ? x5 : ~x1)) | (x6 & ~x7 & ~x1 & x5))) | (x5 & x6 & ~x7 & x1 & x4))) | ((~x3 | (x3 & x5 & x6 & ~x7)) & ((x1 & ~x4) | (x0 & (~x1 | (x1 & x4))))) | (x0 & ~x1 & x3 & (x6 ? ~x5 : x4)))) | (x0 & (((x1 | (~x1 & ~x4 & ~x6)) & (x3 ? ~x5 : ~x2)) | (x5 & ((~x1 & ~x2 & ((x4 & (~x6 | (x6 & ~x7))) | (~x3 & x6 & x7))) | (x1 & x3 & x4 & ~x6))) | (~x1 & ~x2 & ~x4 & x6 & ~x7))) | (x3 & ((~x2 & ((~x0 & ~x5) | (x6 & ~x7 & x1 & x5))) | (x5 & ((~x0 & ((x4 & ~x6) | (~x1 & x6 & ~x7))) | (x7 & (~x4 | (x4 & x6))))))) | (~x0 & ~x2 & ~x3);
  assign z35 = (x0 & (x1 ? (x3 ? (x2 ? (~x4 | (x4 & ~x5)) : x4) : x2) : (x2 | (~x2 & x4 & ~x5)))) | ((x2 ? ~x0 : x1) & (~x3 | (x3 & ~x4))) | (x3 & x4 & ((~x0 & (~x2 | (x2 & ~x5))) | (x1 & x2 & x5))) | (~x1 & ~x2 & ~x4);
  assign z36 = x2 ? ((x4 & (((~x5 | (x5 & (~x6 | (x6 & x7)))) & (x1 ? x3 : ~x0)) | (x3 & x5 & x6 & ~x7 & (~x0 | (x0 & x1))))) | (x0 & (~x1 | (x1 & x3 & ~x4))) | (~x0 & ((x3 & ~x4) | (~x1 & ~x3 & ((x5 & x6 & ~x7) | (~x4 & (~x6 | (x6 & x7))))))) | (x1 & ~x3)) : (~x0 | (x0 & (x1 | (~x1 & (~x4 | (x4 & x5))))));
  assign z37 = x3 ? (((~x6 | (x6 & x7)) & (((~x0 | (x0 & x1)) & (~x4 | (x4 & x5))) | (x0 & ~x1 & (x2 | (~x2 & ~x5))))) | (~x0 & (x5 ? (x6 & ~x7) : x4)) | (x0 & ((x1 & ((x4 & ~x5) | (x6 & ~x7 & ~x2 & x5))) | (x6 & ~x7 & ((x2 & x5) | (~x1 & x4 & ~x5)))))) : (~x0 | (x0 & (~x1 | (x1 & x2))));
  assign z38 = (~x0 & ((x4 & (((~x5 | (x5 & (~x6 | (x6 & x7)))) & (x1 ? x3 : ~x2)) | (x5 & x6 & ~x7 & ~x2 & x3))) | (x3 & ~x4) | (~x3 & (x2 | (~x1 & ~x2 & ((x5 & x6 & ~x7) | (~x4 & (~x6 | (x6 & x7))))))))) | (x0 & ((x3 & ((~x2 & (x1 | (~x1 & ~x4 & x6))) | (x2 & ((x4 & ((x5 & ~x6) | (x1 & (~x5 | (x5 & x6 & x7))))) | (~x1 & (~x5 | (x5 & x6))))) | (~x1 & ~x4 & x5 & ~x6))) | (x2 & (x4 ? ~x3 : x1)) | (~x1 & ~x3 & ~x4))) | (x1 & ((~x2 & ~x3) | (x5 & x6 & ~x7 & x2 & x3 & x4)));
  assign z39 = (x3 & ((~x4 & ((x0 & x2 & ~x5) | (x5 & x7))) | (x0 & ((x2 & ((x5 & x6 & ~x7) | (~x1 & x4 & ~x6))) | (~x5 & (x1 ? ~x2 : (x6 ? x4 : ~x2))) | (x1 & x5 & ((x4 & ~x6) | (~x2 & x6 & ~x7))))) | (~x0 & ~x5) | (x5 & ((~x0 & (x6 ? ~x7 : x4)) | (x4 & x6 & x7))))) | (x0 & ((x1 & (x2 ? (x4 & ~x5) : ~x3)) | ((~x4 | (x4 & x5)) & ((x2 & ~x3) | (x6 & ~x7 & ~x1 & ~x2))) | (~x1 & ((x4 & ((~x3 & ~x5) | (~x2 & x5 & ~x6))) | (~x2 & ~x3 & ((x5 & x6 & x7) | (~x4 & ~x6))))))) | (~x0 & ~x3);
  assign z40 = (x0 & ((x4 & ((~x1 & (~x5 | (x6 & ~x7 & x2 & x5))) | (x3 & ((x1 & ~x2) | (x6 & x7 & x2 & x5))) | (x2 & ((x5 & ~x6) | (x1 & (~x5 | (~x3 & x5 & x6 & ~x7))))))) | (~x4 & ((~x1 & ~x2 & (x6 | (x5 & ~x6))) | (x2 & ~x3 & (~x6 | (x6 & ~x7))))) | (x2 & ~x3 & x5 & x6 & x7))) | (~x0 & ((x3 & (((~x5 | (x5 & (~x6 | (x6 & x7)))) & (x1 ? x4 : ~x2)) | (x5 & x6 & ~x7 & ~x2 & x4))) | (x2 & ~x3) | (~x1 & ~x2 & ~x4 & ((x5 & x6 & ~x7) | (~x3 & (~x6 | (x6 & x7))))))) | (x3 & ((x1 & ((~x2 & ~x4) | (x5 & x6 & ~x7 & x2 & x4))) | (x2 & ~x4))) | (x1 & ~x2 & ~x3);
  assign z41 = ~x0 | (x0 & ((x1 & (~x2 ^ ~x3)) | (~x1 & (~x3 | (~x2 & x3 & ~x5))) | (x2 & x3)));
  assign z42 = ((~x5 | (x5 & x6 & ~x7)) & (~x0 | (x0 & ((x2 & ~x3) | (x1 & (~x2 | (x2 & x3 & ~x4))))))) | (x0 & ((x4 & ((x1 & ((~x5 & ~x6 & x2 & x3) | (x6 & x7 & ~x2 & x5))) | (x6 & (x2 ? ((x5 & x7) | (x3 & (~x5 | (x5 & ~x7)))) : ~x1)))) | (~x1 & ((~x5 & ~x6) | (~x4 & x6 & ~x7)) & (~x2 | (x2 & x3))))) | (x5 & (x4 ? (~x6 | (~x0 & x6 & x7)) : x7));
  assign z43 = (x2 & (x0 ? (((x6 ? x4 : ~x5) & (~x1 | (x1 & ~x3))) | (x5 & ((x4 & ~x6) | (x1 & ((~x4 & x7) | (x3 & x6 & (~x4 ^ x7)))))) | (x1 & ((x3 & ~x5) | (~x3 & ~x4 & x6 & ~x7)))) : (((~x3 | (x3 & ~x4)) & (~x5 | (x5 & x6 & ~x7))) | (x4 & (x3 ? x1 : (x5 & (~x6 | (x6 & x7))))) | (~x4 & x5 & x7)))) | (~x2 & ((x6 & ((~x3 & ((~x0 & ~x1 & ~x4 & x7) | (x1 & x5 & ~x7))) | (x5 & ((x1 & ((x4 & x7) | (x3 & ~x4 & ~x7))) | (~x0 & ((~x1 & (x7 ? x3 : ~x4)) | (x3 & x4 & ~x7))))) | (~x0 & ~x1 & x3 & ~x5))) | (~x6 & ((x4 & ((x1 & x5) | (~x0 & ~x1 & x3))) | (~x0 & ~x1 & ~x4 & (~x5 | (x5 & x7))))) | (x1 & (~x5 | (~x4 & x5 & x7))))) | (x0 & ((~x1 & ~x4 & (x7 ? x5 : x6)) | (x5 & x6 & ~x7 & x1 & x3 & x4)));
  assign z44 = ((x2 ? x3 : ~x1) & (x0 ? (x4 & (~x5 | (x5 & x6))) : ~x4)) | (x3 & (~x1 | (x1 & x2)) & (x0 ? (~x4 | (x4 & x5 & ~x6)) : x4)) | (x2 & ~x3) | (~x2 & (x1 | (x0 & ~x1 & ~x3 & (x6 ? ~x4 : x5))));
  assign z45 = (x0 & (x1 ^ ~x2)) | (~x0 & ((~x4 & (x1 ? (x2 & (x6 | (x5 & ~x6))) : (~x2 & (~x6 | (x6 & ~x7))))) | (~x1 & ~x2 & (x5 ? ((x6 & x7) | (x4 & (~x6 | (x6 & ~x7)))) : x4)))) | (x1 & ~x2) | (~x1 & x2);
  assign z46 = ~x1 | (x1 & ((~x3 & (x2 | (~x4 & x6 & ~x7 & ~x0 & ~x2))) | (x3 & ((x4 & (x5 ? (((~x6 | (x6 & x7)) & (~x0 | (x0 & x2))) | (x2 & x6 & ~x7)) : x2)) | (x2 & ~x4) | (~x0 & ~x2 & (~x5 | (x5 & x6 & ~x7))))) | (~x2 & (x0 | (~x0 & ~x4 & x5 & (~x6 | (x6 & x7)))))));
  assign z47 = ((~x5 | (x5 & (~x6 | (x6 & ~x7)))) & ((x0 & x1 & x2 & x3) | (~x0 & ~x1 & ~x2 & x4))) | (~x0 & ((~x4 & (x1 ? (x2 & (x6 | (x5 & ~x6))) : (~x2 & (~x6 | (x6 & ~x7))))) | (x5 & x6 & x7 & ~x1 & ~x2))) | (~x1 & (x2 | (x0 & ~x2))) | (x1 & (~x2 | (x0 & x2 & (~x3 | (x3 & x4 & x5 & x6 & x7)))));
  assign z48 = (~x3 & (x1 ? x2 : ~x0)) | (x3 & ((x2 & (((x5 ? (x6 & x7) : ~x6) & (x1 ? x4 : ~x0)) | (x1 & ~x4) | (x4 & (~x0 | (x0 & x1)) & (x5 ? (~x6 | (x6 & ~x7)) : x6)))) | (~x0 & ~x1 & ~x4 & (x5 ? (~x6 | (x6 & ~x7)) : x6)))) | (x0 & ~x1) | (x1 & ~x2);
  assign z49 = ((~x0 | (x0 & x1)) & (~x2 | (x2 & x3 & x4))) | (x0 & ~x1) | (x2 & ((x1 & ~x3) | (~x4 & ((x1 & x3) | (~x0 & ~x1 & (x6 | (x5 & ~x6)))))));
  assign z50 = (x4 & (((~x5 | (x5 & (~x6 | (x6 & ~x7)))) & (x0 ? (x1 & x3) : ~x2)) | (x3 & x5 & x6 & x7 & x0 & x1 & x2))) | (x2 & (~x0 | (x3 & ~x4 & x0 & x1))) | (~x2 & ((x5 & x6 & x7) | (~x4 & (~x6 | (x6 & ~x7)))) & (~x0 | (x0 & x1 & x3))) | (x0 & (~x1 | (x1 & ~x3)));
  assign z51 = x0 ? (~x1 | (x1 & ((~x2 & ((x6 & (((~x5 | (x5 & ~x7)) & (~x4 | (x3 & x4))) | (x3 & x5 & x7))) | (x3 & ~x6 & (~x5 | (x4 & x5))))) | (~x4 & (x6 ? x2 : x5))))) : ((~x3 & (~x1 | (x1 & x2))) | (x1 & (~x2 | (x2 & x3 & ~x4))) | (x3 & ((~x1 & ~x4 & (x6 | (x5 & ~x6))) | (x2 & x4))));
  assign z52 = (x3 & ((x0 & (((~x5 | (x5 & x6)) & (x1 ? (~x2 | (x2 & ~x4)) : x2)) | (x4 & x5 & ~x6 & (x2 | (x1 & ~x2))))) | (x5 & ((x4 & x6 & x1 & x2) | (~x0 & ~x1 & ~x4 & ~x6))) | (~x0 & (x1 ? (~x2 | (x2 & ~x4)) : (x4 ? x2 : x6))) | (x4 & ~x5 & x1 & x2))) | (~x1 & ((x0 & ~x2) | (x2 & ~x3 & ~x4 & x6))) | (~x2 & ((~x0 & ~x3) | (x0 & x1 & ~x4 & x5 & ~x6))) | (~x4 & ((x0 & ((x1 & ~x3 & x6) | (x2 & x5 & ~x6))) | (~x0 & x2 & ~x3 & x5 & ~x6))) | (~x0 & x1 & x2 & ((x4 & x5 & ~x6) | (~x3 & (~x5 | (x5 & x6)))));
  assign z53 = (x5 & (((~x6 | (x6 & ~x7)) & ((~x1 & ((x3 & x4) | (x0 & ~x2 & ~x3))) | (x1 & ((x0 & ((~x3 & x4) | (x2 & x3 & ~x4))) | (~x0 & x2 & x3 & x4))) | (~x0 & (x2 ? (x3 & ~x4) : ~x3)))) | (x6 & ((x7 & ((x4 & (x2 ? (x0 ? (~x1 ^ ~x3) : x3) : (~x1 | (x1 & ~x3)))) | (~x0 & x1 & x2 & x3 & ~x4))) | (x0 & x1 & x2 & ~x3 & ~x4))) | (x1 & ~x4 & ~x6 & (~x2 ^ ~x3)))) | (~x5 & ((~x1 & ((x3 & x4) | (x0 & ~x2 & ~x3))) | (~x0 & (x2 ? (x3 & ~x4) : ~x3)) | (x1 & ((x2 & (x0 ? (~x4 & (~x3 | (x3 & x6))) : (x3 & x4))) | (x0 & ~x3 & x4))))) | (~x4 & ((x0 & (x1 ? (~x2 & ~x3) : (x2 & x3))) | (x1 & x6 & ((~x2 & x3) | (~x0 & x2 & ~x3))) | (~x1 & ~x2 & x3))) | (~x1 & x2 & ~x3);
  assign z54 = (x5 & ((x3 & ((~x1 & ((~x0 & ((~x2 & ~x6) | (x4 & x6 & x7))) | (x2 & x4 & (~x6 | (x6 & ~x7))))) | (x1 & ((x4 & ((x0 & (x6 ? ~x7 : x2)) | (~x2 & (~x6 | (x6 & x7))))) | (x2 & ~x4 & (~x6 | (x6 & (~x7 | (x0 & x7))))))) | (x6 & ((x0 & x2 & x4 & x7) | (~x0 & ~x2 & ~x7))))) | (~x3 & (x0 ? x1 : x2) & (~x6 | (x6 & (~x7 | (x4 & x7))))) | (~x0 & x1 & ~x2 & ~x4 & ~x6))) | (~x2 & ((~x0 & ((x3 & ~x5) | (~x4 & x6 & x1 & ~x3))) | (x0 & x3 & (~x1 | (x1 & (~x4 | (x4 & ~x5))))) | (~x1 & ~x3))) | (x2 & (x3 ? ((~x1 & ~x4) | (~x5 & (x1 ? ((~x4 & x6) | (x0 & (~x6 | (x4 & x6)))) : x4))) : (x0 ? ~x1 : ~x5))) | (x0 & x1 & ~x3 & ~x5);
  assign z55 = ~x1 | (x1 & ((~x4 & (x0 ? (x3 & (x6 ? ~x2 : x5)) : (x6 | (x5 & ~x6)))) | (x0 & ((~x3 & (~x2 | (x2 & x5 & ~x6))) | (x2 & (~x5 | (x5 & ((x6 & ~x7) | (x4 & (x6 ? x7 : x3))))))))));
  assign z56 = (x3 & ((x2 & (((~x4 | (x0 & x4)) & (~x1 | (x1 & (~x5 | (x5 & x6 & ~x7))))) | (x5 & ((~x0 & x4 & (~x6 | (x6 & ~x7))) | (x0 & x1 & ~x4 & x6 & x7))) | (~x0 & x4 & ~x5))) | (x1 & ((~x4 & ((x6 & x7 & ~x2 & x5) | (~x0 & ((x5 & ~x6) | (~x2 & x6 & ~x7))))) | (x0 & ((~x2 & (~x5 | (x5 & x6 & ~x7))) | (x5 & (~x6 | (x4 & x6 & x7))))))))) | (~x2 & (~x1 | (x1 & ~x3))) | (x2 & (x0 ? ~x3 : (x5 ? ((x4 & x6 & x7) | (~x3 & (~x6 | (x6 & ~x7)))) : ~x3)));
  assign z57 = (x2 & ((x3 & ((~x1 & (x0 | (~x0 & x5 & ~x6))) | (x5 & ((x6 & (x0 ? (x1 & (~x4 ^ x7)) : (~x7 | (x4 & x7)))) | (x1 & ~x4 & ~x6))) | (~x5 & (~x0 | (x0 & x1 & ~x4))))) | (~x1 & ~x3) | (x1 & (((~x5 | (x5 & (~x6 | (x6 & ~x7)))) & (x0 ? x4 : ~x3)) | (~x3 & ((x0 & ~x4) | (x4 & x5 & x6 & x7))))))) | (~x1 & ~x2) | (x1 & ((~x2 & ((~x3 & (x0 | (x6 & ~x7 & ~x0 & ~x4))) | (~x0 & ~x4 & x5 & (~x6 | (x6 & x7))) | (x3 & (x0 ? (~x4 & (x6 ? ~x7 : x5)) : (~x5 | (x5 & x6 & (~x7 | (x4 & x7)))))))) | (x3 & x5 & ((~x0 & x4 & ~x6) | (x6 & x7 & x0 & ~x4)))));
  assign z58 = (~x1 & ((x0 & (~x2 | (x2 & ~x3))) | (~x0 & ~x3) | (x3 & ((x2 & (~x4 | (x4 & x5 & x6 & x7))) | (~x0 & (((~x6 | (x6 & ~x7)) & (x4 ? x5 : ~x2)) | (x4 & ~x5) | (x6 & x7 & ~x2 & x5))))))) | (x1 & ~x2) | (x2 & (x3 ? ((x0 & (((~x5 | (x5 & x6 & ~x7)) & (x4 | (x1 & ~x4))) | (x4 & x5 & (~x6 | (x1 & x6 & x7))))) | (x1 & ~x4 & (x6 ? ~x0 : x5))) : x1));
  assign z59 = (x1 & ((x0 & (x3 ? ((~x5 & (x2 ^ x4)) | (x5 & ((x6 & (x2 ? (~x4 | (x4 & x7)) : (x7 | (x4 & ~x7)))) | (~x2 & x4 & ~x6))) | (~x2 & ~x4 & (~x6 | (x6 & ~x7)))) : (~x2 | (x2 & ~x4 & (x6 | (x5 & ~x6)))))) | (~x0 & x2 & ~x3) | (x4 & (~x5 | (x5 & (~x6 | (x6 & ~x7)))) & (x2 ? x3 : ~x0)))) | (~x0 & ((x2 & ((x3 & (~x4 | (x4 & x5 & x6 & x7))) | (~x1 & ~x3 & ((x5 & x6 & x7) | (~x4 & (~x6 | (x6 & ~x7))))))) | ((~x6 | (x6 & ~x7)) & ((~x2 & ~x4) | (~x1 & x4 & x5))) | (~x1 & x4 & ~x5) | (x6 & x7 & ~x2 & x5))) | (x0 & (x2 ? ((~x1 & (~x3 | (x3 & ~x4 & x6))) | (x3 & ~x4 & x5 & ~x6)) : ~x1));
  assign z60 = (~x0 & ((x5 & (((~x6 | (x6 & ~x7)) & ((x2 & x3 & ~x4) | (~x1 & (x3 ? x4 : ~x2)))) | (x4 & x6 & x7 & (x2 ? x3 : ~x1)))) | (~x5 & ((x2 & x3 & ~x4) | (~x1 & (x3 ? x4 : ~x2)))) | (x2 & ~x3) | (~x2 & (x3 ? ~x4 : x1)))) | (x0 & ~x1) | (x1 & (x2 ? ((x3 & (((~x5 | (x5 & (~x6 | (x6 & ~x7)))) & (x4 | (x0 & ~x4))) | (x5 & x6 & x7 & (~x4 | (x0 & x4))))) | (x0 & ~x3 & ~x4)) : (x4 ? x3 : x0)));
  assign z61 = ~x0 | (x0 & (~x2 | (x2 & (~x3 | (x3 & ((~x4 & (x6 ? ~x1 : x5)) | (x1 & (~x5 | (x5 & (x6 | (x4 & ~x6)))))))))));
  assign z62 = ~x0 | (x0 & (~x1 | (x1 & ((~x4 & (x6 ? ~x3 : x5)) | (x3 & (~x5 | (x5 & (x6 | (x4 & ~x6)))))))));
endmodule