module pla__e64 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55,
    x56, x57, x58, x59, x60, x61, x62, x63, x64,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54,
    x55, x56, x57, x58, x59, x60, x61, x62, x63, x64;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64;
  assign z00 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x47 & ~x46 & x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x00 & ~x03;
  assign z01 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & x05 & ~x04 & ~x00 & ~x03;
  assign z02 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x44 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x38 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x32 & ~x31 & ~x30 & x29 & ~x28 & x27 & ~x26 & ~x25 & ~x24 & ~x23 & ~x22 & ~x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z03 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & x44 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x38 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x32 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x23 & ~x22 & ~x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z04 = x15 & x29;
  assign z05 = x29;
  assign z06 = ~x43 & ~x37 & x29 & ~x28 & x14 & ~x15;
  assign z07 = x43 & ~x37 & x29 & ~x15 & ~x28;
  assign z08 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & x38 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x32 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x23 & ~x22 & ~x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z09 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x32 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & x23 & ~x22 & ~x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z10 = ~x37 & x29 & ~x15 & x28;
  assign z11 = x37 & ~x15 & x29;
  assign z12 = ~x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x03 & x06;
  assign z13 = ~x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & x41 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x03 & ~x07;
  assign z14 = ~x58 & x50 & ~x43 & ~x37 & x29 & ~x28 & ~x15 & ~x10 & ~x14;
  assign z15 = ~x58 & ~x43 & ~x37 & x29 & ~x28 & ~x15 & x10 & ~x14;
  assign z16 = ~x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & x26 & ~x25 & ~x24 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x03 & ~x07;
  assign z17 = ~x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & x03 & ~x07;
  assign z18 = x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x11 & ~x10 & ~x07 & ~x08;
  assign z19 = x64 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z20 = ~x62 & ~x60 & ~x58 & ~x56 & x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & ~x00 & ~x03;
  assign z21 = ~x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & x00 & ~x03;
  assign z22 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & x36 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z23 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x21 & ~x18 & ~x17 & x16 & ~x15 & ~x14 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z24 = ~x60 & ~x58 & ~x50 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x10 & x11;
  assign z25 = ~x60 & ~x58 & ~x50 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & x29 & ~x28 & ~x25 & x24 & ~x15 & ~x10 & ~x14;
  assign z26 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & x32 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x21 & ~x20 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z27 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x21 & ~x20 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z28 = ~x60 & ~x58 & ~x50 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & x29 & ~x28 & x25 & ~x15 & ~x10 & ~x14;
  assign z29 = x60 & ~x58 & ~x50 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & x29 & ~x28 & ~x15 & ~x10 & ~x14;
  assign z30 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x21 & ~x18 & ~x17 & ~x15 & ~x14 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z31 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & x21 & ~x18 & ~x17 & ~x15 & ~x14 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z32 = ~x58 & ~x50 & x46 & ~x43 & ~x40 & ~x39 & ~x37 & x29 & ~x28 & ~x15 & ~x10 & ~x14;
  assign z33 = ~x58 & ~x50 & ~x43 & ~x40 & x39 & ~x37 & x29 & ~x28 & ~x15 & ~x10 & ~x14;
  assign z34 = x58 & ~x43 & ~x37 & x29 & ~x28 & ~x14 & ~x15;
  assign z35 = ~x62 & ~x61 & ~x60 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & x04 & ~x00 & ~x03;
  assign z36 = ~x62 & x61 & ~x60 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & ~x00 & ~x03;
  assign z37 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x32 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x21 & ~x20 & x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z38 = ~x62 & ~x61 & ~x60 & x59 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z39 = ~x62 & ~x61 & ~x60 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z40 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & x54 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z41 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & x33 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z42 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & x49 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z43 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & x01;
  assign z44 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x00 & x02;
  assign z45 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & x34 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z46 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & x09 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z47 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z48 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z49 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & x53 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x04 & ~x00 & ~x03;
  assign z50 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z51 = ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x49 & x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z52 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z53 = ~x64 & x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x17 & ~x15 & ~x14 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z54 = ~x62 & ~x60 & ~x58 & ~x56 & x55 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & ~x00 & ~x03;
  assign z55 = ~x62 & ~x60 & ~x58 & ~x56 & ~x51 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & x35 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x06 & ~x00 & ~x03;
  assign z56 = ~x64 & ~x63 & ~x62 & ~x61 & ~x60 & ~x59 & ~x58 & ~x57 & ~x56 & ~x55 & ~x54 & ~x53 & ~x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x47 & ~x46 & ~x45 & ~x43 & ~x42 & ~x41 & ~x40 & ~x39 & ~x37 & ~x36 & ~x35 & ~x34 & ~x33 & ~x31 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & ~x21 & x20 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x07 & ~x06 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z57 = ~x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & ~x22 & x18 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x03 & ~x06;
  assign z58 = ~x62 & ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x41 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x26 & ~x25 & ~x24 & x22 & ~x15 & ~x14 & ~x11 & ~x10 & ~x08 & ~x07 & ~x03 & ~x06;
  assign z59 = ~x58 & ~x50 & ~x43 & x40 & ~x37 & x29 & ~x28 & ~x15 & ~x10 & ~x14;
  assign z60 = ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x11 & ~x10 & x07 & ~x08;
  assign z61 = ~x60 & ~x58 & ~x56 & ~x50 & ~x47 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x11 & x08 & ~x10;
  assign z62 = ~x60 & ~x58 & ~x56 & ~x50 & x47 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x10 & ~x11;
  assign z63 = ~x60 & ~x58 & x56 & ~x50 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & ~x30 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x10 & ~x11;
  assign z64 = ~x60 & ~x58 & ~x50 & ~x46 & ~x43 & ~x40 & ~x39 & ~x37 & x30 & x29 & ~x28 & ~x25 & ~x24 & ~x15 & ~x14 & ~x10 & ~x11;
endmodule