module pla__ex4 ( 
    x000, x001, x002, x003, x004, x005, x006, x007, x008, x009, x010, x011,
    x012, x013, x014, x015, x016, x017, x018, x019, x020, x021, x022, x023,
    x024, x025, x026, x027, x028, x029, x030, x031, x032, x033, x034, x035,
    x036, x037, x038, x039, x040, x041, x042, x043, x044, x045, x046, x047,
    x048, x049, x050, x051, x052, x053, x054, x055, x056, x057, x058, x059,
    x060, x061, x062, x063, x064, x065, x066, x067, x068, x069, x070, x071,
    x072, x073, x074, x075, x076, x077, x078, x079, x080, x081, x082, x083,
    x084, x085, x086, x087, x088, x089, x090, x091, x092, x093, x094, x095,
    x096, x097, x098, x099, x100, x101, x102, x103, x104, x105, x106, x107,
    x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119,
    x120, x121, x122, x123, x124, x125, x126, x127,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27  );
  input  x000, x001, x002, x003, x004, x005, x006, x007, x008, x009,
    x010, x011, x012, x013, x014, x015, x016, x017, x018, x019, x020, x021,
    x022, x023, x024, x025, x026, x027, x028, x029, x030, x031, x032, x033,
    x034, x035, x036, x037, x038, x039, x040, x041, x042, x043, x044, x045,
    x046, x047, x048, x049, x050, x051, x052, x053, x054, x055, x056, x057,
    x058, x059, x060, x061, x062, x063, x064, x065, x066, x067, x068, x069,
    x070, x071, x072, x073, x074, x075, x076, x077, x078, x079, x080, x081,
    x082, x083, x084, x085, x086, x087, x088, x089, x090, x091, x092, x093,
    x094, x095, x096, x097, x098, x099, x100, x101, x102, x103, x104, x105,
    x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117,
    x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27;
  assign z00 = x040 & ((~x000 & ~x080 & (x032 | x072) & (x008 | x048)) | (~x016 & ~x064 & (x048 | x072) & (x008 | x032)) | (~x032 & ~x048) | (~x008 & ~x072));
  assign z01 = x041 & ((~x001 & ~x081 & (x033 | x073) & (x009 | x049)) | (~x017 & ~x065 & (x049 | x073) & (x009 | x033)) | (~x033 & ~x049) | (~x009 & ~x073));
  assign z02 = x042 & ((~x002 & ~x082 & (x034 | x074) & (x010 | x050)) | (~x018 & ~x066 & (x050 | x074) & (x010 | x034)) | (~x034 & ~x050) | (~x010 & ~x074));
  assign z03 = x043 & ((~x003 & ~x083 & (x035 | x075) & (x011 | x051)) | (~x019 & ~x067 & (x051 | x075) & (x011 | x035)) | (~x035 & ~x051) | (~x011 & ~x075));
  assign z04 = x044 & ((~x004 & ~x084 & (x036 | x076) & (x012 | x052)) | (~x020 & ~x068 & (x052 | x076) & (x012 | x036)) | (~x036 & ~x052) | (~x012 & ~x076));
  assign z05 = x045 & ((x053 & ((x077 & (x085 ? (((~x109 | ~x117) & ((~x005 & (x037 | x069) & (x013 | x021 | x061 | x093)) | (~x029 & (x013 | x021) & (x061 | x093)) | ~x013 | ~x021)) | ((x061 | x093) & (((~x101 | ~x125) & ((~x005 & (x037 | x069)) | (~x029 & (x013 | x021)))) | (~x029 & (x013 | x021) & (~x005 | ~x037 | ~x069)))) | ((~x061 | ~x093) & (~x037 | ~x069 | (~x005 & (x013 | x021) & (x037 | x069 | x109 | x117)))) | (~x005 & (((x037 | x069) & (x013 | x021) & (~x029 | ~x101 | ~x125)) | ((x109 | x117) & (x013 | x021) & (~x029 | ~x125))))) : ~x005)) | (~x021 & ~x069 & (x013 | x037)) | (~x005 & x037 & ~x085))) | (x013 & ((~x005 & ~x085 & (x037 | x077)) | (~x021 & ~x069 & x077))) | (~x037 & ~x053) | (~x069 & x077 & ~x021 & x037) | (~x013 & ~x077));
  assign z06 = x046 & ((x054 & ((x078 & (x086 ? (((~x110 | ~x118) & ((~x006 & (x038 | x070) & (x014 | x022 | x062 | x094)) | (~x030 & (x014 | x022) & (x062 | x094)) | ~x014 | ~x022)) | ((x062 | x094) & (((~x102 | ~x126) & ((~x006 & (x038 | x070)) | (~x030 & (x014 | x022)))) | (~x030 & (x014 | x022) & (~x006 | ~x038 | ~x070)))) | ((~x062 | ~x094) & (~x038 | ~x070 | (~x006 & (x014 | x022) & (x038 | x070 | x110 | x118)))) | (~x006 & (((x038 | x070) & (x014 | x022) & (~x030 | ~x102 | ~x126)) | ((x110 | x118) & (x014 | x022) & (~x030 | ~x126))))) : ~x006)) | (~x022 & ~x070 & (x014 | x038)) | (~x006 & x038 & ~x086))) | (x014 & ((~x006 & ~x086 & (x038 | x078)) | (~x022 & ~x070 & x078))) | (~x038 & ~x054) | (~x070 & x078 & ~x022 & x038) | (~x014 & ~x078));
  assign z08 = ~x040 & ((~x048 & ((~x072 & (x080 ? x000 : (((x104 | x112) & ((x000 & (~x032 | ~x064) & (~x008 | ~x016 | ~x056 | ~x088)) | (x024 & (~x008 | ~x016) & (~x056 | ~x088)) | x008 | x016)) | ((~x056 | ~x088) & ((x024 & (~x008 | ~x016) & (x000 | x032 | x064 | x096 | x120)) | (x000 & (~x032 | ~x064) & (x096 | x120)))) | ((x056 | x088) & ((x000 & (~x008 | ~x016) & (~x032 | ~x064 | ~x104 | ~x112)) | x032 | x064)) | (x000 & (((~x032 | ~x064) & (~x008 | ~x016) & (x024 | x096 | x120)) | ((~x104 | ~x112) & (~x008 | ~x016) & (x024 | x120))))))) | (x016 & x064 & (~x008 | ~x032)) | (x000 & ~x032 & x080))) | (~x008 & ((x000 & x080 & (~x032 | ~x072)) | (x016 & x064 & ~x072))) | (x032 & x048) | (x064 & ~x072 & x016 & ~x032) | (x008 & x072));
  assign z09 = ~x041 & ((x001 & x081 & (~x033 | ~x073) & (~x009 | ~x049)) | (x017 & x065 & (~x049 | ~x073) & (~x009 | ~x033)) | (x033 & x049) | (x009 & x073));
  assign z10 = ~x042 & ((x002 & x082 & (~x034 | ~x074) & (~x010 | ~x050)) | (x018 & x066 & (~x050 | ~x074) & (~x010 | ~x034)) | (x034 & x050) | (x010 & x074));
  assign z11 = ~x043 & ((x003 & x083 & (~x035 | ~x075) & (~x011 | ~x051)) | (x019 & x067 & (~x051 | ~x075) & (~x011 | ~x035)) | (x035 & x051) | (x011 & x075));
  assign z12 = ~x044 & ((x004 & x084 & (~x036 | ~x076) & (~x012 | ~x052)) | (x020 & x068 & (~x052 | ~x076) & (~x012 | ~x036)) | (x036 & x052) | (x012 & x076));
  assign z13 = ~x045 & ((~x053 & ((~x077 & (x085 ? x005 : (((x109 | x117) & ((x005 & (~x037 | ~x069) & (~x013 | ~x021 | ~x061 | ~x093)) | x013 | x021 | (x029 & (~x013 | ~x021) & (~x061 | ~x093)))) | ((~x061 | ~x093) & ((x029 & (~x013 | ~x021) & (x005 | x037 | x069 | x101 | x125)) | (x005 & (~x037 | ~x069) & (x101 | x125)))) | ((x061 | x093) & (x037 | x069 | (x005 & (~x013 | ~x021) & (~x109 | ~x117 | ~x037 | ~x069)))) | (x005 & (((~x037 | ~x069) & (~x013 | ~x021) & (x029 | x101 | x125)) | ((~x109 | ~x117) & (~x013 | ~x021) & (x029 | x125))))))) | (x021 & x069 & (~x013 | ~x037)) | (x005 & ~x037 & x085))) | (~x013 & ((x005 & x085 & (~x037 | ~x077)) | (x021 & x069 & ~x077))) | (x037 & x053) | (x069 & ~x077 & x021 & ~x037) | (x013 & x077));
  assign z14 = ~x046 & ((~x054 & ((~x078 & (x086 ? x006 : (((x110 | x118) & ((x006 & (~x038 | ~x070) & (~x014 | ~x022 | ~x062 | ~x094)) | x014 | x022 | (x030 & (~x014 | ~x022) & (~x062 | ~x094)))) | ((~x062 | ~x094) & ((x030 & (~x014 | ~x022) & (x006 | x038 | x070 | x102 | x126)) | (x006 & (~x038 | ~x070) & (x102 | x126)))) | ((x062 | x094) & (x038 | x070 | (x006 & (~x014 | ~x022) & (~x110 | ~x118 | ~x038 | ~x070)))) | (x006 & (((~x038 | ~x070) & (~x014 | ~x022) & (x030 | x102 | x126)) | ((~x110 | ~x118) & (~x014 | ~x022) & (x030 | x126))))))) | (x022 & x070 & (~x014 | ~x038)) | (x006 & ~x038 & x086))) | (~x014 & ((x006 & x086 & (~x038 | ~x078)) | (x022 & x070 & ~x078))) | (x038 & x054) | (x070 & ~x078 & x022 & ~x038) | (x014 & x078));
  assign z07 = 1'b0;
  assign z15 = 1'b0;
  assign z16 = 1'b0;
  assign z17 = 1'b0;
  assign z18 = 1'b0;
  assign z19 = 1'b0;
  assign z20 = 1'b0;
  assign z21 = 1'b0;
  assign z22 = 1'b0;
  assign z23 = 1'b0;
  assign z24 = 1'b0;
  assign z25 = 1'b0;
  assign z26 = 1'b0;
  assign z27 = 1'b0;
endmodule