module pla__misex3c ( 
    di__larrow__11__rarrow__, di__larrow__10__rarrow__,
    di__larrow__9__rarrow__, di__larrow__8__rarrow__,
    di__larrow__7__rarrow__, di__larrow__6__rarrow__,
    di__larrow__5__rarrow__, di__larrow__4__rarrow__,
    di__larrow__3__rarrow__, di__larrow__2__rarrow__,
    di__larrow__1__rarrow__, di__larrow__0__rarrow__,
    ci__larrow__1__rarrow__, ci__larrow__0__rarrow__,
    d__larrow__7__rarrow__, d__larrow__6__rarrow__, d__larrow__5__rarrow__,
    d__larrow__4__rarrow__, d__larrow__3__rarrow__, d__larrow__2__rarrow__,
    d__larrow__1__rarrow__, d__larrow__0__rarrow__,
    cd__larrow__1__rarrow__, cd__larrow__0__rarrow__,
    c__larrow__1__rarrow__, c__larrow__0__rarrow__,
    cs__larrow__0__rarrow__, v__larrow__0__rarrow__  );
  input  di__larrow__11__rarrow__, di__larrow__10__rarrow__,
    di__larrow__9__rarrow__, di__larrow__8__rarrow__,
    di__larrow__7__rarrow__, di__larrow__6__rarrow__,
    di__larrow__5__rarrow__, di__larrow__4__rarrow__,
    di__larrow__3__rarrow__, di__larrow__2__rarrow__,
    di__larrow__1__rarrow__, di__larrow__0__rarrow__,
    ci__larrow__1__rarrow__, ci__larrow__0__rarrow__;
  output d__larrow__7__rarrow__, d__larrow__6__rarrow__,
    d__larrow__5__rarrow__, d__larrow__4__rarrow__, d__larrow__3__rarrow__,
    d__larrow__2__rarrow__, d__larrow__1__rarrow__, d__larrow__0__rarrow__,
    cd__larrow__1__rarrow__, cd__larrow__0__rarrow__,
    c__larrow__1__rarrow__, c__larrow__0__rarrow__,
    cs__larrow__0__rarrow__, v__larrow__0__rarrow__;
  assign d__larrow__7__rarrow__ = (di__larrow__9__rarrow__ & (di__larrow__7__rarrow__ ? (~di__larrow__6__rarrow__ & ci__larrow__0__rarrow__) : (~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__))) | (~di__larrow__6__rarrow__ & ((di__larrow__10__rarrow__ & ~di__larrow__8__rarrow__ & ~di__larrow__7__rarrow__) | (~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__ & di__larrow__8__rarrow__ & di__larrow__7__rarrow__))) | (di__larrow__10__rarrow__ & ((~di__larrow__8__rarrow__ & di__larrow__7__rarrow__ & (ci__larrow__1__rarrow__ | (di__larrow__6__rarrow__ & di__larrow__5__rarrow__))) | (~di__larrow__7__rarrow__ & ((ci__larrow__0__rarrow__ & (~di__larrow__5__rarrow__ | (di__larrow__6__rarrow__ & di__larrow__5__rarrow__))) | (di__larrow__8__rarrow__ & ci__larrow__1__rarrow__))))) | (di__larrow__8__rarrow__ & ((~di__larrow__11__rarrow__ & ci__larrow__1__rarrow__) | (~di__larrow__9__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & ci__larrow__0__rarrow__))) | (~di__larrow__8__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & ~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__);
  assign d__larrow__6__rarrow__ = (ci__larrow__0__rarrow__ & ((di__larrow__9__rarrow__ & (di__larrow__7__rarrow__ ^ di__larrow__6__rarrow__)) | (~di__larrow__10__rarrow__ & di__larrow__7__rarrow__))) | (ci__larrow__1__rarrow__ & ((~di__larrow__10__rarrow__ & (~di__larrow__7__rarrow__ | (di__larrow__8__rarrow__ & di__larrow__7__rarrow__))) | (di__larrow__8__rarrow__ & (~di__larrow__11__rarrow__ | (di__larrow__10__rarrow__ & ~di__larrow__7__rarrow__) | (di__larrow__11__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__))))) | (~ci__larrow__0__rarrow__ & ((di__larrow__8__rarrow__ & (di__larrow__7__rarrow__ ? (~di__larrow__6__rarrow__ & ~ci__larrow__1__rarrow__) : di__larrow__6__rarrow__)) | (~di__larrow__9__rarrow__ & di__larrow__7__rarrow__ & ~ci__larrow__1__rarrow__)));
  assign d__larrow__5__rarrow__ = (di__larrow__7__rarrow__ & ((~di__larrow__10__rarrow__ & (ci__larrow__0__rarrow__ | (di__larrow__6__rarrow__ & ci__larrow__1__rarrow__))) | (~di__larrow__9__rarrow__ & ((~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__) | (di__larrow__8__rarrow__ & di__larrow__6__rarrow__ & ci__larrow__0__rarrow__))) | (~di__larrow__6__rarrow__ & ~ci__larrow__1__rarrow__) | (~di__larrow__8__rarrow__ & di__larrow__6__rarrow__ & ((~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__) | (di__larrow__10__rarrow__ & di__larrow__5__rarrow__))))) | (di__larrow__10__rarrow__ & ((di__larrow__6__rarrow__ & ci__larrow__1__rarrow__ & di__larrow__11__rarrow__ & ~di__larrow__8__rarrow__) | (di__larrow__8__rarrow__ & ~di__larrow__6__rarrow__ & ci__larrow__0__rarrow__))) | (di__larrow__6__rarrow__ & ci__larrow__1__rarrow__ & (~di__larrow__11__rarrow__ | (di__larrow__8__rarrow__ & ~di__larrow__7__rarrow__)));
  assign d__larrow__4__rarrow__ = (di__larrow__10__rarrow__ & ~di__larrow__7__rarrow__ & (di__larrow__6__rarrow__ ? (di__larrow__5__rarrow__ & ci__larrow__0__rarrow__) : ~di__larrow__8__rarrow__)) | (di__larrow__5__rarrow__ & (ci__larrow__0__rarrow__ ? (~di__larrow__10__rarrow__ | (di__larrow__7__rarrow__ & (~di__larrow__9__rarrow__ | ~di__larrow__6__rarrow__))) : ~ci__larrow__1__rarrow__)) | (di__larrow__3__rarrow__ & ci__larrow__1__rarrow__);
  assign d__larrow__3__rarrow__ = ci__larrow__1__rarrow__ ? ((di__larrow__4__rarrow__ & ~di__larrow__1__rarrow__ & (di__larrow__2__rarrow__ | (di__larrow__5__rarrow__ & di__larrow__0__rarrow__))) | (di__larrow__1__rarrow__ & (~di__larrow__4__rarrow__ | (di__larrow__5__rarrow__ & (~di__larrow__2__rarrow__ | (di__larrow__2__rarrow__ & di__larrow__0__rarrow__)))))) : (di__larrow__3__rarrow__ ? (di__larrow__2__rarrow__ ? ~di__larrow__1__rarrow__ : di__larrow__4__rarrow__) : di__larrow__1__rarrow__);
  assign d__larrow__2__rarrow__ = ci__larrow__1__rarrow__ ? ((di__larrow__4__rarrow__ & (~di__larrow__2__rarrow__ ^ ~di__larrow__1__rarrow__)) | (~di__larrow__5__rarrow__ & di__larrow__2__rarrow__)) : ((di__larrow__3__rarrow__ & (di__larrow__2__rarrow__ ? ~di__larrow__1__rarrow__ : di__larrow__4__rarrow__)) | (~di__larrow__4__rarrow__ & di__larrow__1__rarrow__));
  assign d__larrow__1__rarrow__ = (ci__larrow__1__rarrow__ & ((di__larrow__5__rarrow__ & ((di__larrow__3__rarrow__ & ~di__larrow__1__rarrow__) | (di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__))) | (di__larrow__2__rarrow__ & (~di__larrow__5__rarrow__ | (di__larrow__4__rarrow__ & ~di__larrow__1__rarrow__))))) | (di__larrow__2__rarrow__ & (~di__larrow__4__rarrow__ | (~ci__larrow__1__rarrow__ & (~di__larrow__3__rarrow__ | (di__larrow__3__rarrow__ & ~di__larrow__1__rarrow__)))));
  assign d__larrow__0__rarrow__ = di__larrow__0__rarrow__ & (~di__larrow__5__rarrow__ | (~di__larrow__4__rarrow__ & di__larrow__2__rarrow__) | (~di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | ~ci__larrow__1__rarrow__ | (di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & ~di__larrow__1__rarrow__ & ci__larrow__1__rarrow__));
  assign cd__larrow__1__rarrow__ = di__larrow__9__rarrow__ ? ci__larrow__1__rarrow__ : (~di__larrow__8__rarrow__ & ~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__ & ((di__larrow__0__rarrow__ & ((di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ((~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | (di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__))) | (~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__))) | (~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__1__rarrow__ & ~di__larrow__0__rarrow__)));
  assign cd__larrow__0__rarrow__ = (~ci__larrow__1__rarrow__ & (di__larrow__5__rarrow__ ? ((di__larrow__7__rarrow__ & ((di__larrow__0__rarrow__ & ((~di__larrow__9__rarrow__ & ~ci__larrow__0__rarrow__ & ((di__larrow__8__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | (~di__larrow__8__rarrow__ & di__larrow__6__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__))) | (~di__larrow__10__rarrow__ & di__larrow__9__rarrow__ & di__larrow__8__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & ci__larrow__0__rarrow__))) | (di__larrow__9__rarrow__ & di__larrow__8__rarrow__ & di__larrow__6__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ~di__larrow__0__rarrow__ & (di__larrow__10__rarrow__ | ~ci__larrow__0__rarrow__)))) | (di__larrow__9__rarrow__ & di__larrow__8__rarrow__ & ~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & di__larrow__0__rarrow__ & ~ci__larrow__0__rarrow__ & ((~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | (di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__)))) : ((di__larrow__8__rarrow__ & di__larrow__6__rarrow__) | (~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__0__rarrow__)))) | (di__larrow__8__rarrow__ & ((di__larrow__10__rarrow__ & ((~di__larrow__6__rarrow__ & ci__larrow__0__rarrow__) | (~di__larrow__7__rarrow__ & ci__larrow__1__rarrow__))) | (~di__larrow__10__rarrow__ & ((di__larrow__6__rarrow__ & ci__larrow__0__rarrow__) | (di__larrow__7__rarrow__ & ci__larrow__1__rarrow__))) | (di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & ((di__larrow__11__rarrow__ & ci__larrow__1__rarrow__) | (~di__larrow__9__rarrow__ & ci__larrow__0__rarrow__))) | (~di__larrow__7__rarrow__ & di__larrow__5__rarrow__ & ci__larrow__0__rarrow__))) | (~di__larrow__8__rarrow__ & ((di__larrow__11__rarrow__ & ci__larrow__1__rarrow__ & (di__larrow__7__rarrow__ | (di__larrow__10__rarrow__ & di__larrow__6__rarrow__))) | (~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & di__larrow__0__rarrow__)));
  assign c__larrow__1__rarrow__ = (di__larrow__8__rarrow__ & ((~di__larrow__11__rarrow__ & ci__larrow__1__rarrow__) | (di__larrow__5__rarrow__ & ((~di__larrow__6__rarrow__ & di__larrow__0__rarrow__ & ~ci__larrow__1__rarrow__ & ((di__larrow__3__rarrow__ & ~di__larrow__1__rarrow__ & ((di__larrow__7__rarrow__ & (~di__larrow__4__rarrow__ ^ ~di__larrow__2__rarrow__) & ((~di__larrow__10__rarrow__ & di__larrow__9__rarrow__ & ci__larrow__0__rarrow__) | (~di__larrow__9__rarrow__ & ~ci__larrow__0__rarrow__))) | (di__larrow__9__rarrow__ & ~di__larrow__7__rarrow__ & di__larrow__4__rarrow__ & ~di__larrow__2__rarrow__ & ~ci__larrow__0__rarrow__))) | (di__larrow__9__rarrow__ & ~di__larrow__7__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__))) | (~di__larrow__7__rarrow__ & ci__larrow__0__rarrow__))))) | (~di__larrow__8__rarrow__ & di__larrow__0__rarrow__ & ((~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__) | (~di__larrow__9__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & ~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__))) | (~di__larrow__2__rarrow__ & ~di__larrow__0__rarrow__);
  assign c__larrow__0__rarrow__ = (di__larrow__0__rarrow__ & ((di__larrow__5__rarrow__ & (ci__larrow__1__rarrow__ ? (di__larrow__1__rarrow__ ? di__larrow__2__rarrow__ : di__larrow__4__rarrow__) : ((di__larrow__8__rarrow__ & (di__larrow__9__rarrow__ ? ((di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & (((di__larrow__10__rarrow__ | ~ci__larrow__0__rarrow__) & ((di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | (~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__))) | (~di__larrow__10__rarrow__ & di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ci__larrow__0__rarrow__))) | (~di__larrow__10__rarrow__ & di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__4__rarrow__ & di__larrow__1__rarrow__ & ci__larrow__0__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__)) : (di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~ci__larrow__0__rarrow__ & ((~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | (di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__))))) | (di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & ~di__larrow__9__rarrow__ & ~di__larrow__8__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__)))) | (~di__larrow__8__rarrow__ & di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__))) | (~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & ~di__larrow__0__rarrow__ & ~ci__larrow__1__rarrow__);
  assign cs__larrow__0__rarrow__ = (di__larrow__0__rarrow__ & (di__larrow__8__rarrow__ ? (di__larrow__9__rarrow__ ? ((di__larrow__4__rarrow__ & ((di__larrow__3__rarrow__ & ((di__larrow__10__rarrow__ & ((di__larrow__6__rarrow__ & ((~ci__larrow__0__rarrow__ & ((~di__larrow__11__rarrow__ & ~di__larrow__7__rarrow__ & ~di__larrow__1__rarrow__ & ci__larrow__1__rarrow__ & (di__larrow__5__rarrow__ ^ di__larrow__2__rarrow__)) | (di__larrow__11__rarrow__ & di__larrow__7__rarrow__ & di__larrow__5__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__))) | (di__larrow__7__rarrow__ & di__larrow__5__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & ~ci__larrow__1__rarrow__))) | (~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ~ci__larrow__1__rarrow__))) | (di__larrow__5__rarrow__ & ~ci__larrow__1__rarrow__ & ((di__larrow__7__rarrow__ & ((~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ci__larrow__0__rarrow__ & ~di__larrow__10__rarrow__ & ~di__larrow__6__rarrow__) | (di__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__ & di__larrow__6__rarrow__ & di__larrow__2__rarrow__))) | (~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__))))) | (~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ~ci__larrow__1__rarrow__ & (~di__larrow__10__rarrow__ | ~ci__larrow__0__rarrow__)))) | (~di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ~di__larrow__4__rarrow__ & di__larrow__2__rarrow__ & ~ci__larrow__1__rarrow__ & ((~di__larrow__10__rarrow__ & di__larrow__7__rarrow__ & ci__larrow__0__rarrow__ & (di__larrow__3__rarrow__ ^ di__larrow__1__rarrow__)) | (~di__larrow__7__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__1__rarrow__ & (di__larrow__10__rarrow__ | ~ci__larrow__0__rarrow__))))) : (di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ~ci__larrow__1__rarrow__ & ~ci__larrow__0__rarrow__ & ((di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__) | (~di__larrow__4__rarrow__ & di__larrow__2__rarrow__ & (di__larrow__3__rarrow__ ^ di__larrow__1__rarrow__))))) : (~ci__larrow__0__rarrow__ & ((~di__larrow__9__rarrow__ & ~ci__larrow__1__rarrow__ & ((di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ((~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | (di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__))) | (~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__))) | (~di__larrow__11__rarrow__ & di__larrow__10__rarrow__ & di__larrow__9__rarrow__ & ~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & ci__larrow__1__rarrow__))))) | (~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__1__rarrow__ & ~di__larrow__0__rarrow__ & ~ci__larrow__1__rarrow__ & ((di__larrow__9__rarrow__ & di__larrow__8__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & di__larrow__2__rarrow__ & (di__larrow__10__rarrow__ | ~ci__larrow__0__rarrow__)) | (~di__larrow__9__rarrow__ & ~di__larrow__8__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & ~ci__larrow__0__rarrow__)));
  assign v__larrow__0__rarrow__ = (~ci__larrow__0__rarrow__ & ((ci__larrow__1__rarrow__ & ((di__larrow__8__rarrow__ & ((~di__larrow__9__rarrow__ & ((~di__larrow__10__rarrow__ & di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__) | (~di__larrow__11__rarrow__ & ~di__larrow__7__rarrow__))) | (~di__larrow__5__rarrow__ & ((di__larrow__11__rarrow__ & di__larrow__10__rarrow__ & di__larrow__9__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__) | (~di__larrow__11__rarrow__ & ~di__larrow__7__rarrow__ & ~di__larrow__2__rarrow__))) | ((~di__larrow__4__rarrow__ | ~di__larrow__3__rarrow__) & ((~di__larrow__11__rarrow__ & ~di__larrow__7__rarrow__) | (di__larrow__11__rarrow__ & di__larrow__10__rarrow__ & di__larrow__9__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__))) | (~di__larrow__11__rarrow__ & ~di__larrow__7__rarrow__ & (di__larrow__1__rarrow__ | (di__larrow__5__rarrow__ & di__larrow__2__rarrow__))) | (di__larrow__11__rarrow__ & di__larrow__10__rarrow__ & di__larrow__9__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & (~di__larrow__2__rarrow__ | ~di__larrow__1__rarrow__ | ~di__larrow__0__rarrow__)))) | (~di__larrow__7__rarrow__ & ((di__larrow__9__rarrow__ & ((~di__larrow__10__rarrow__ & ~di__larrow__6__rarrow__) | (di__larrow__11__rarrow__ & di__larrow__10__rarrow__ & ~di__larrow__8__rarrow__))) | (~di__larrow__6__rarrow__ & ((~di__larrow__8__rarrow__ & (di__larrow__3__rarrow__ | di__larrow__2__rarrow__ | ~di__larrow__0__rarrow__)) | (~di__larrow__11__rarrow__ & ~di__larrow__1__rarrow__))))) | (~di__larrow__1__rarrow__ & (((di__larrow__11__rarrow__ | di__larrow__7__rarrow__) & ((~di__larrow__5__rarrow__ & di__larrow__2__rarrow__) | (di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__))) | (~di__larrow__2__rarrow__ & ~di__larrow__0__rarrow__) | (~di__larrow__5__rarrow__ & (~di__larrow__0__rarrow__ | (~di__larrow__8__rarrow__ & di__larrow__2__rarrow__))))) | (~di__larrow__11__rarrow__ & (~di__larrow__10__rarrow__ | (di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__ & di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__))) | (~di__larrow__5__rarrow__ & ~di__larrow__4__rarrow__) | (~di__larrow__10__rarrow__ & ((di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__ & di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__) | (~di__larrow__9__rarrow__ & ~di__larrow__8__rarrow__ & di__larrow__6__rarrow__))))) | (~ci__larrow__1__rarrow__ & (di__larrow__9__rarrow__ ? ((di__larrow__3__rarrow__ & ((di__larrow__8__rarrow__ & di__larrow__7__rarrow__ & di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ~di__larrow__4__rarrow__) | (~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & di__larrow__1__rarrow__))) | (di__larrow__2__rarrow__ & ((~di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & di__larrow__4__rarrow__) | (~di__larrow__4__rarrow__ & ~di__larrow__1__rarrow__ & di__larrow__0__rarrow__))) | (~di__larrow__6__rarrow__ & (di__larrow__7__rarrow__ ? (~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__) : ((di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__) | (~di__larrow__4__rarrow__ & ~di__larrow__2__rarrow__)))) | (di__larrow__7__rarrow__ & ((~di__larrow__2__rarrow__ & ((di__larrow__4__rarrow__ & ~di__larrow__1__rarrow__) | (di__larrow__8__rarrow__ & di__larrow__6__rarrow__ & di__larrow__5__rarrow__))) | (di__larrow__8__rarrow__ & di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ((di__larrow__4__rarrow__ & (~di__larrow__1__rarrow__ | ~di__larrow__0__rarrow__)) | (~di__larrow__3__rarrow__ & di__larrow__0__rarrow__)))))) : ((~di__larrow__4__rarrow__ & ((~di__larrow__8__rarrow__ & di__larrow__3__rarrow__) | (di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ~di__larrow__2__rarrow__))) | (di__larrow__4__rarrow__ & ((di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & (~di__larrow__3__rarrow__ | (di__larrow__5__rarrow__ & di__larrow__2__rarrow__))) | (~di__larrow__8__rarrow__ & (~di__larrow__3__rarrow__ | ~di__larrow__0__rarrow__ | (~di__larrow__5__rarrow__ & ~di__larrow__1__rarrow__))))) | (~di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & (~di__larrow__8__rarrow__ | (di__larrow__7__rarrow__ & di__larrow__3__rarrow__ & di__larrow__1__rarrow__))) | (~di__larrow__8__rarrow__ & ((~di__larrow__2__rarrow__ & di__larrow__1__rarrow__) | (di__larrow__6__rarrow__ & di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__)))))) | (di__larrow__0__rarrow__ & ((~di__larrow__9__rarrow__ & ((~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__) | (di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__))) | (di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & (~di__larrow__8__rarrow__ | ~di__larrow__7__rarrow__ | ~di__larrow__6__rarrow__)) | (~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__2__rarrow__ & (di__larrow__8__rarrow__ | di__larrow__7__rarrow__ | di__larrow__6__rarrow__)))) | (~di__larrow__8__rarrow__ & ~di__larrow__7__rarrow__ & di__larrow__4__rarrow__ & ~di__larrow__2__rarrow__ & (~di__larrow__6__rarrow__ | (di__larrow__5__rarrow__ & di__larrow__3__rarrow__ & ~di__larrow__1__rarrow__))) | (~di__larrow__4__rarrow__ & ~di__larrow__0__rarrow__ & (di__larrow__3__rarrow__ ? ~di__larrow__1__rarrow__ : (di__larrow__2__rarrow__ & di__larrow__1__rarrow__))))) | (~ci__larrow__1__rarrow__ & ((di__larrow__9__rarrow__ & ((~di__larrow__8__rarrow__ & (di__larrow__4__rarrow__ ? (~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__) : ~di__larrow__3__rarrow__)) | (di__larrow__4__rarrow__ & ((di__larrow__10__rarrow__ & di__larrow__8__rarrow__ & (di__larrow__7__rarrow__ ? (di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & (~di__larrow__1__rarrow__ | ~di__larrow__0__rarrow__)) : (~di__larrow__6__rarrow__ & (di__larrow__2__rarrow__ | (~di__larrow__3__rarrow__ & ci__larrow__0__rarrow__))))) | (di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__ & ~di__larrow__5__rarrow__ & di__larrow__3__rarrow__))) | (di__larrow__10__rarrow__ & di__larrow__8__rarrow__ & (di__larrow__7__rarrow__ ? (di__larrow__6__rarrow__ & di__larrow__5__rarrow__ & ((~di__larrow__4__rarrow__ & di__larrow__3__rarrow__) | ~di__larrow__2__rarrow__ | (~di__larrow__3__rarrow__ & di__larrow__0__rarrow__))) : (~di__larrow__6__rarrow__ & ((~di__larrow__4__rarrow__ & ~di__larrow__2__rarrow__) | (di__larrow__3__rarrow__ & di__larrow__1__rarrow__))))) | (~di__larrow__6__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__0__rarrow__))) | ((di__larrow__4__rarrow__ ? (~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__) : (~di__larrow__3__rarrow__ & di__larrow__1__rarrow__)) & ((di__larrow__8__rarrow__ & di__larrow__6__rarrow__) | (di__larrow__10__rarrow__ & di__larrow__7__rarrow__ & ci__larrow__0__rarrow__))) | (~di__larrow__9__rarrow__ & ((~di__larrow__8__rarrow__ & (di__larrow__7__rarrow__ ? (di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__) : di__larrow__5__rarrow__)) | (~di__larrow__7__rarrow__ & (di__larrow__4__rarrow__ ? (~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__) : (~di__larrow__3__rarrow__ & di__larrow__0__rarrow__))) | (di__larrow__5__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__1__rarrow__) | (di__larrow__8__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__) | (~di__larrow__10__rarrow__ & ci__larrow__0__rarrow__) | (di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__ & di__larrow__6__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__))) | (ci__larrow__0__rarrow__ & ((di__larrow__2__rarrow__ & ((di__larrow__4__rarrow__ & ((~di__larrow__10__rarrow__ & ((di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__) | (di__larrow__3__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__))) | (di__larrow__3__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__ & (~di__larrow__8__rarrow__ | ~di__larrow__6__rarrow__)))) | (~di__larrow__6__rarrow__ & ((~di__larrow__7__rarrow__ & ~di__larrow__5__rarrow__) | (di__larrow__10__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__1__rarrow__))) | (~di__larrow__8__rarrow__ & ~di__larrow__4__rarrow__ & ~di__larrow__1__rarrow__))) | (~di__larrow__10__rarrow__ & ((~di__larrow__7__rarrow__ & ((~di__larrow__4__rarrow__ & ~di__larrow__3__rarrow__) | (di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__))) | (~di__larrow__4__rarrow__ & ((~di__larrow__1__rarrow__ & ~di__larrow__0__rarrow__) | (di__larrow__7__rarrow__ & ~di__larrow__6__rarrow__ & ~di__larrow__2__rarrow__))) | (~di__larrow__6__rarrow__ & ((~di__larrow__5__rarrow__ & di__larrow__3__rarrow__) | (di__larrow__7__rarrow__ & (di__larrow__3__rarrow__ ? di__larrow__1__rarrow__ : di__larrow__4__rarrow__)))))) | (~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ~di__larrow__0__rarrow__))) | (~di__larrow__4__rarrow__ & ((~di__larrow__7__rarrow__ & ((di__larrow__3__rarrow__ & di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__) | (di__larrow__5__rarrow__ & ~di__larrow__3__rarrow__ & ~di__larrow__0__rarrow__))) | (di__larrow__6__rarrow__ & (di__larrow__3__rarrow__ ? (di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__) : ~di__larrow__5__rarrow__)) | (~di__larrow__3__rarrow__ & di__larrow__0__rarrow__ & (~di__larrow__5__rarrow__ | ~di__larrow__1__rarrow__)))) | (~di__larrow__7__rarrow__ & ((di__larrow__2__rarrow__ & di__larrow__1__rarrow__ & di__larrow__0__rarrow__ & di__larrow__5__rarrow__ & di__larrow__4__rarrow__ & di__larrow__3__rarrow__) | (~di__larrow__6__rarrow__ & ~di__larrow__5__rarrow__ & (di__larrow__3__rarrow__ ? ~di__larrow__2__rarrow__ : di__larrow__1__rarrow__)))) | (di__larrow__4__rarrow__ & ~di__larrow__2__rarrow__ & ~di__larrow__1__rarrow__ & ~di__larrow__0__rarrow__)));
endmodule