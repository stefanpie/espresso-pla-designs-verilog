module pla__Z9sym ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z0;
  assign z0 = (~x4 & (x3 ? ((~x2 & (x1 ? ((x0 & (~x5 | (x5 & x6 & ~x7))) | (x5 & (~x6 | (x6 & x7 & ~x8))) | (~x0 & ((~x5 & (x8 ? ~x6 : x7)) | (x6 & (~x7 | (x7 & x8)))))) : ((x8 & (x0 ? (x6 ? x7 : ~x5) : ((x5 & ~x6) | (x6 & ~x7) | (~x5 & x7)))) | (x0 & ((x6 & ~x7) | (~x5 & x7 & ~x8))) | (x7 & ~x8 & ~x0 & x6)))) | (~x0 & ((x2 & (x5 ? (x6 ? (~x7 ^ ~x8) : (~x7 | (x7 & x8))) : ((x6 & (~x7 | (x7 & x8))) | (~x1 & (x8 ? ~x6 : x7))))) | (~x1 & x5 & (x6 ? (~x7 ^ x8) : (x7 & ~x8))))) | (x2 & ((x0 & ((~x7 & (x1 ? (~x5 ^ ~x6) : (x5 & x6))) | (~x1 & ~x5))) | (x1 & ((~x5 & ~x6) | (~x8 & (x5 ? (~x6 ^ ~x7) : (x6 & x7))))))) | (x0 & ~x1 & x5 & (~x6 | (x6 & x7 & ~x8)))) : ((x0 & ((x5 & ((x6 & ~x7 & x1 & x2) | (~x6 & x8 & ~x1 & ~x2))) | (((~x5 & (x8 ? ~x6 : x7)) | (x6 & (~x7 | (x7 & x8)))) & (x1 ^ x2)) | (~x5 & ((x1 & x2) | (x7 & x8 & ~x1 & ~x2))) | (~x1 & ~x2 & x6 & (~x7 ^ ~x8)))) | (~x0 & (((x1 ^ x2) & ((x6 & (~x7 ^ ~x8)) | (x8 & (x5 ? ~x6 : x7)))) | (x1 & x2 & ((~x5 & (x8 ? ~x6 : x7)) | (x6 & (~x7 | (x7 & x8))))) | (~x1 & ~x2 & x6 & x7 & x8))) | (x1 & x2 & x5 & (~x6 | (x6 & x7 & ~x8)))))) | (~x3 & ((x4 & (x5 ? ((x2 & (x7 ? ((~x0 & (x6 ^ x8)) | (x1 & ~x6 & ~x8)) : ((x0 & (x1 ^ x6)) | (~x0 & (~x6 | (x6 & x8))) | (x1 & x6 & ~x8)))) | (x0 & x1 & ~x2 & x6 & ~x7)) : (x2 ? ((x0 & (~x1 | (x1 & x6 & ~x7))) | (x1 & (~x6 | (x6 & x7 & ~x8))) | (~x0 & ((x6 & (~x7 | (x7 & x8))) | (~x1 & (x8 ? ~x6 : x7))))) : (((x8 ? ~x6 : x7) & (x0 ^ x1)) | (x0 & x1) | (x7 & x8 & ~x0 & ~x1))))) | (x5 & (((x1 ? (~x2 & ~x8) : (x2 ^ x8)) & (x0 ? (x6 & x7) : (~x6 ^ ~x7))) | ((x1 ^ x2) & ((x0 & ~x6) | (x7 & x8 & ~x0 & x6))) | (~x1 & ~x2 & ~x8 & (x0 ? (~x6 ^ ~x7) : (x6 & x7))))))) | (x4 & (((~x5 ^ ~x6) & ((~x0 & ((~x2 & (x1 ? (~x7 | (x7 & x8)) : (~x7 ^ ~x8))) | (x3 & ((~x1 & (~x7 ^ x8)) | (x2 & (~x7 ^ ~x8)))))) | (x3 & ((x0 & (x1 ? (~x2 & ~x7) : (x7 ? ~x8 : x2))) | (x1 & ~x8 & (~x2 ^ ~x7)))) | (x0 & ~x1 & ~x2 & (~x7 | (x7 & x8))))) | (x5 & x6 & (((~x7 ^ ~x8) & (x0 ? (~x1 & ~x2) : (x1 ? ~x2 : x3))) | (~x0 & ((~x1 & ~x2 & (~x7 ^ x8)) | (~x7 & ~x8 & x2 & x3))) | (x3 & ~x7 & ~x8 & (x1 ? ~x2 : x0)))) | (x3 & ~x5 & ~x6 & ((x0 & (~x1 | (x1 & x2 & ~x7))) | (x1 & (~x2 | (x2 & x7 & ~x8))) | (~x0 & ((~x1 & (x8 ? ~x2 : x7)) | (x2 & (~x7 | (x7 & x8)))))))));
endmodule