module pla__duke2 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28;
  assign z00 = ~x09 & ~x18 & ((x17 & (x05 ? (~x07 | ~x15) : (x07 ? x15 : (~x15 | (~x00 & x15))))) | (x04 & ~x05 & ~x07 & x12 & ~x14 & ~x15 & ~x17 & ~x21));
  assign z01 = ~x17 & ((~x05 & ((~x07 & x18 & ((~x09 & ((~x15 & ((x06 & ~x08 & (~x21 | (~x14 & x21)) & (x02 ^ x11)) | (~x02 & x08 & x11 & x13 & ~x14 & ~x21 & (~x10 | (x04 & x10 & ~x12))))) | (~x02 & x08 & x11 & x15 & ~x21))) | (~x02 & x08 & x09 & x11 & x15))) | (x02 & x07 & ~x09 & x11 & x15 & ~x18))) | (~x04 & x05 & ~x07 & x08 & ~x09 & ~x11 & x15 & x18 & ~x21));
  assign z02 = ~x17 & ((~x09 & ((~x05 & ((x01 & x07 & ~x15 & ~x18 & (x08 | x16)) | (x18 & ((~x07 & ((x06 & (~x02 | ~x11)) | (~x08 & x15))) | (x08 & x15 & x21))))) | (x18 & ((~x07 & ((~x04 & ((~x06 & ~x15) | (x05 & x08 & ~x11 & x15 & ~x21))) | (x05 & (x08 ? (x15 & x21) : ~x15)) | (~x06 & ~x12 & ~x15))) | (x05 & x08 & ~x15 & x21))))) | (x08 & x18 & ((~x07 & (((x09 | ~x21) & ((x02 & ~x05 & ~x11 & x15) | (~x04 & x05 & x12 & ~x15))) | (~x05 & ~x15))) | (x05 & ~x15 & (x07 | ~x12)) | (~x05 & x15 & (~x02 | x07)))));
  assign z03 = (~x09 & (x05 ? ((~x07 & ((x17 & ~x18) | (~x08 & ~x15 & ~x17 & x18))) | (x07 & x08 & ~x15 & ~x17 & x18)) : ((x07 & x08 & x15 & ~x17 & x18) | (x17 & ~x18)))) | (~x05 & ~x07 & x08 & ~x17 & x18 & x09 & ~x15);
  assign z04 = ~x14 & ~x20;
  assign z05 = ~x05 & ~x07 & ~x09 & ~x14 & ~x15 & ~x17 & x18 & ((x02 & ((x06 & ~x08 & ~x11 & x21) | (~x06 & x08 & ~x10 & x13 & ~x21))) | (x06 & ((~x02 & ~x08 & x11 & x21) | (x08 & x10 & x12 & ~x13 & x16 & ~x21))) | (~x06 & ((~x08 & x21 & (x04 ^ x12)) | (x08 & x10 & x12 & ~x13 & ~x16 & ~x21))));
  assign z06 = ~x09 & ((~x05 & ((~x07 & ((~x17 & x18 & ((~x02 & x08 & x11 & x15 & ~x21) | (~x15 & ((~x14 & ((x06 & ((~x02 & ~x08 & x11 & x21) | (x08 & x10 & x12 & ~x13 & x16 & ~x21))) | (x08 & ~x21 & (((~x10 | (x04 & x10 & ~x12)) & (~x13 | (~x02 & x11 & x13))) | (~x06 & ((x02 & ~x10 & x13) | (x10 & x12 & ~x13 & ~x16))))) | (x04 & ~x06 & ~x08 & ~x12 & x21))) | (~x08 & ~x21 & ((~x02 & x06 & x11) | (x04 & ~x06 & ~x12))))))) | (x17 & ~x18 & x00 & x15))) | (x17 & ~x18 & x07 & ~x15))) | (~x07 & x08 & x04 & x05 & ~x12 & ~x15 & ~x17 & x18 & ~x21));
  assign z07 = ~x17 & x18 & ((~x09 & (~x07 ^ x08) & (x05 ^ x15)) | (~x05 & ~x07 & x08 & x09 & ~x15 & x16));
  assign z08 = x14 & ~x20;
  assign z09 = (~x17 & ((x18 & ((~x07 & ((~x15 & ((~x09 & ((~x21 & ((x04 & ~x12 & ((~x05 & ~x06 & ~x08) | (x02 & x08 & x13 & ~x14))) | (~x05 & ((x02 & x08 & x13 & ~x14 & (~x10 | (x10 & x12))) | (~x02 & x06 & ~x08 & x11))))) | (x05 & ~x08 & ~x19))) | (~x04 & x05 & x08 & x12 & (x09 | ~x21)))) | (x08 & x15 & ((x02 & ~x05 & ~x11 & (x09 | ~x21)) | (x05 & ~x09 & x21))))) | (x05 & x08 & ~x15 & (x07 | ~x12 | (~x09 & x21))))) | (x04 & ~x05 & ~x07 & ~x09 & x12 & ~x14 & ~x15 & ~x18 & ~x21))) | (~x07 & ~x09 & ~x15 & x17 & ~x18);
  assign z10 = (~x07 & ((~x09 & ((x05 & ((x17 & ~x18) | (~x15 & ~x17 & x18 & ~x06 & ~x08))) | (x15 & ~x17 & x18 & ~x05 & ~x06 & ~x08))) | (~x15 & ~x17 & x18 & ~x05 & x08 & x09))) | (~x15 & ~x17 & x18 & x05 & x07 & x08) | (x17 & ~x18 & ~x05 & ~x09);
  assign z11 = ~x18 & ~x17 & ~x15 & ~x09 & x07 & x01 & ~x05;
  assign z12 = ~x09 & ((~x07 & ((~x17 & x18 & ~x21 & ((~x04 & ((x05 & x08 & ~x11 & x15) | (~x05 & ~x06 & ~x08 & x12 & ~x15))) | (~x05 & ((~x15 & (x08 ? (~x14 & (~x10 | (x04 & x10 & ~x12)) & (~x13 | (~x02 & x11 & x13))) : ((x04 & ~x06 & ~x12) | (x06 & (x02 ^ x11))))) | (~x02 & x08 & x11 & x15))) | (x04 & x05 & x08 & ~x12 & ~x15))) | (x00 & ~x05 & x15 & x17 & ~x18))) | (~x15 & x17 & ~x18 & ~x05 & x07));
  assign z13 = ~x09 & x17 & ~x18 & (~x05 | (x05 & ~x07));
  assign z14 = (~x17 & ((x08 & x18 & (x07 ? (~x19 & (x05 ^ x15)) : ((x09 | (~x09 & ~x21)) & ((x11 & x15 & ~x02 & ~x05) | (~x12 & ~x15 & x04 & x05))))) | (~x05 & ~x09 & ~x18 & ((x07 & x15 & (~x02 | ~x11 | (x02 & x11))) | (x04 & ~x07 & x12 & ~x14 & ~x15 & ~x21))))) | (~x05 & ~x09 & ~x18 & (x07 ? (~x01 | x17) : (x15 & x17)));
  assign z15 = ~x18 & x17 & ~x15 & ~x09 & x05 & ~x07;
  assign z16 = x08 & ~x17 & x18 & (x05 ? (x09 & ~x15 & (x07 | ~x12)) : ((~x07 & ~x15 & (x09 ? ~x19 : (~x14 & ~x21 & ((x06 & ((x02 & ((x04 & ~x12) | (~x10 & x13))) | (x12 & ~x16 & ((~x02 & x11) | (x10 & ~x13))))) | ((~x10 | (x04 & x10 & ~x12)) & (~x13 | (~x02 & x11 & x13))) | (~x06 & x12 & x16 & ((~x02 & x11) | (x10 & ~x13))))))) | (x09 & x15 & (~x02 | x07))));
  assign z17 = ~x09 & ((~x05 & ((x17 & ~x18 & x07 & ~x15) | (~x07 & ((x17 & ~x18 & x00 & x15) | (~x08 & ~x15 & ~x17 & x18 & (~x21 | (~x14 & x21)) & ((x02 & x06 & ~x11) | (~x04 & ~x06 & x12))))))) | (~x04 & x05 & ~x07 & x08 & ~x11 & x15 & ~x17 & x18 & ~x21));
  assign z18 = ~x05 & ~x07 & ~x09 & ~x17 & x18 & ((~x14 & ~x15 & ((x02 & ((x06 & ~x08 & ~x11 & x21) | (~x06 & x08 & ~x10 & x13 & ~x21))) | (x12 & ((~x06 & ((~x04 & ~x08 & x21) | (~x13 & ~x16 & ~x21 & x08 & x10))) | (~x13 & x16 & ~x21 & x06 & x08 & x10))))) | (~x08 & x15 & x19));
  assign z19 = ~x18 & x17 & ~x15 & ~x09 & ~x05 & ~x07;
  assign z20 = ~x07 & ~x17 & ((~x09 & ((x18 & ((~x21 & (x04 ? (~x12 & ~x15 & (x05 ? x08 : (x08 ? (x10 & ~x14 & (~x13 | (~x02 & x11 & x13))) : ~x06))) : ((x05 & x08 & ~x11 & x15) | (~x05 & ~x06 & ~x08 & x12 & ~x15)))) | (~x05 & ~x06 & ~x08 & ~x14 & ~x15 & x21 & (x04 ^ x12)))) | (x04 & ~x05 & x12 & ~x14 & ~x15 & ~x18 & ~x21))) | (x04 & x05 & x08 & x09 & ~x12 & ~x15 & x18));
  assign z21 = ~x17 & x18 & ((~x07 & ((~x05 & ((~x06 & ~x08 & ~x09 & x15) | (x09 & ~x15 & x06 & x08))) | (x05 & x06 & ~x08 & ~x09 & ~x15))) | (~x05 & x07 & x08 & ~x09 & x15));
  assign z22 = ~x17 & x18 & ((~x07 & ((x05 & x06 & ~x08 & ~x09 & ~x15) | (~x05 & ((x06 & ~x08 & ~x09 & x15) | (x08 & x09 & ~x15))))) | (~x05 & x07 & x08 & x15));
  assign z23 = x18 & ~x17 & ~x15 & x09 & x08 & ~x05 & ~x07;
  assign z24 = ~x09 & ~x17 & ((~x07 & ((~x21 & ((x04 & ~x15 & ((x05 & x08 & ~x12 & x18) | (~x05 & x12 & ~x14 & ~x18))) | (x08 & x15 & x18 & ((~x02 & ~x05 & x11) | (~x04 & x05 & ~x11))))) | (~x15 & x18 & ~x05 & ~x08))) | (x01 & ~x05 & x07 & x08 & ~x15 & ~x18));
  assign z25 = ~x05 & ~x07 & ~x17 & x18 & (x08 ? (x09 & ~x15) : (~x09 & x15));
  assign z26 = ~x20 & (x14 | x21);
  assign z27 = (~x09 & ((~x17 & x18 & (x07 ? (x08 & x19 & (x05 ^ x15)) : ((~x21 & ((~x04 & ((x05 & x08 & ~x11 & x15) | (~x05 & ~x06 & ~x08 & x12 & ~x15))) | (x02 & ~x05 & x06 & ~x08 & ~x11 & ~x15))) | (x05 & ~x08 & ~x15 & x19)))) | (~x05 & x17 & ~x18 & ((x07 & ~x15) | (x00 & ~x07 & x15))))) | (~x07 & x08 & x03 & ~x05 & x09 & ~x15 & ~x17 & x18 & x19);
  assign z28 = (~x17 & ((x18 & ((~x07 & (x05 ? (x08 & ((~x04 & x12 & ~x15 & (x09 | ~x21)) | (~x09 & x15 & x21))) : ((~x09 & ((~x14 & ((~x02 & x11 & ((~x15 & x21 & x06 & ~x08) | (x08 & x10 & x12 & ~x21))) | (~x15 & ((x04 & ~x06 & ~x08 & ~x12 & x21) | (x08 & x10 & x12 & ~x21 & (~x13 | (x02 & x13))))))) | (~x08 & x15 & ~x19))) | (x02 & x08 & ~x11 & x15 & (x09 | ~x21))))) | (~x05 & x08 & x15 & (~x02 | x07 | (~x09 & x21))))) | (~x05 & x07 & ~x09 & x15 & ~x18 & (~x02 | ~x11)))) | (~x09 & x17 & ~x18 & (x05 ? ~x07 : (x15 & (~x07 | ~x19))));
endmodule