module pla__apex4 ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18;
  assign z01 = (x1 & (x2 ? (x4 ? ((~x3 & ((x0 & ~x6 & ~x7 & (x5 | (~x5 & ~x8))) | (~x0 & ~x5 & x6 & x7))) | (x6 & x7 & ~x8 & ~x0 & x3 & x5)) : ((x5 & ((~x3 & ((x0 & ~x7 & (x6 | (~x6 & ~x8))) | (x6 & x7 & ~x8))) | (~x0 & x3 & (x6 ? (~x7 & ~x8) : (x7 & x8))))) | (~x3 & ~x5 & x6 & ((x0 & (~x7 ^ x8)) | (~x7 & x8))))) : (x3 ? (x4 & ((~x0 & ((x7 & x8 & ~x5 & ~x6) | (~x7 & ~x8 & x5 & x6))) | (x6 & x7 & x0 & x5))) : (~x4 & (x5 ? (x7 & ~x8) : (~x7 & x8)) & (x0 ^ x6))))) | (x0 & ((~x2 & ((~x1 & ((x5 & ((~x3 & x4 & x6 & ~x7 & x8) | (x7 & ~x8 & ~x4 & ~x6))) | (x4 & ((~x3 & ~x5 & (x6 ? (~x7 & ~x8) : (x7 & x8))) | (x7 & ~x8 & x3 & ~x6))) | (x3 & ~x4 & (x6 ? x7 : (~x7 & (x8 | (~x5 & ~x8))))))) | (x5 & ~x6 & x8 & (x3 ? (x4 & x7) : (~x4 & ~x7))))) | (~x1 & x3 & ((x2 & ((x6 & ((x5 & (x4 ? x7 : (~x7 ^ x8))) | (x4 & ~x5 & (~x7 ^ ~x8)))) | (x4 & x5 & ~x6 & ~x7))) | (x4 & ~x5 & ~x6 & ~x7 & ~x8))))) | (~x1 & x2 & x3 & x4 & ~x7 & x8 & x5 & x6);
  assign z02 = (x2 & ((x0 & ((~x5 & ((x3 & ((x1 & ((~x7 & x8 & ~x4 & x6) | (x4 & ~x6 & ~x8))) | (~x4 & ((x6 & ~x7 & ~x8) | (~x1 & x7 & (x8 | (x6 & ~x8))))) | (~x7 & ~x8 & ~x1 & ~x6))) | (~x6 & ((~x3 & ((~x1 & (x4 ? (x7 & ~x8) : ~x7)) | (~x7 & ~x8 & x1 & ~x4))) | (x8 & (x4 ^ x7)))) | (~x1 & x6 & ((~x7 & ~x8) | (x7 & x8 & ~x3 & ~x4))))) | (x5 & ((x3 & ((~x1 & ((~x4 & ~x6 & (~x7 ^ ~x8)) | (~x7 & ~x8 & x4 & x6))) | (x1 & ((~x6 & ~x7) | (x4 & x6 & (x7 | (~x7 & x8))))) | (x7 & x8 & ~x4 & ~x6))) | (~x4 & ((~x1 & ((x6 & ~x7 & x8) | (~x3 & ~x6 & x7))) | (x1 & ~x3 & x6 & x7 & x8))) | (~x3 & x4 & x7))) | (~x3 & x7 & x8 & (x1 ? (x4 & x6) : ~x6)))) | (~x0 & ((~x6 & (x7 ? ((x4 & ((x1 & (x5 ? ~x8 : x3)) | (~x5 & x8 & ~x1 & x3))) | (x3 & ~x4 & ~x5)) : (((x5 | (~x5 & ~x8)) & (x1 ? (x3 & ~x4) : (~x3 & x4))) | (x1 & x4 & (x3 ? (~x8 | (~x5 & x8)) : (x5 & x8)))))) | (x6 & (x1 ? ((~x3 & x5 & ((x7 & x8) | (x4 & ~x7 & ~x8))) | (x3 & x4 & ~x5 & x7 & x8)) : ((x3 & (x4 ? (x7 | (~x7 & ~x8)) : (x5 & ~x7))) | (~x3 & ~x4 & x5 & x7 & x8)))) | (x1 & x3 & x4 & x5 & ~x7 & x8))) | (x1 & ~x5 & x8 & ((x3 & ~x6 & (~x4 ^ x7)) | (~x3 & x4 & x6 & ~x7))))) | (~x2 & ((x1 & ((~x5 & (x3 ? ((x4 & ((x6 & ~x7 & x8) | (x0 & x7 & ~x8))) | (x0 & ((~x6 & x7 & x8) | (~x4 & ~x7 & ~x8))) | (x7 & ~x8 & ~x0 & ~x6)) : ((x4 & (x0 ? (x6 & ~x7) : (x8 & (~x6 ^ x7)))) | (~x6 & ~x7 & ~x8) | (x0 & ~x4 & x7 & (x6 ^ ~x8))))) | (x0 & ((~x3 & ((~x7 & ~x8 & x5 & x6) | (x4 & ~x6 & x7))) | (x5 & ((~x6 & ((x3 & ((~x7 & x8) | (x4 & x7 & ~x8))) | (x4 & ~x7 & x8))) | (x7 & ~x8 & x3 & ~x4))))) | (~x0 & x5 & ((~x4 & ((~x7 & (x3 ? (~x6 ^ ~x8) : (~x6 & ~x8))) | (x7 & x8 & ~x3 & x6))) | (x6 & ~x7 & x8 & x3 & x4))))) | (x0 & ((~x1 & ((x3 & ((~x5 & (x4 ? (~x6 & x8) : (x6 ? (~x7 & x8) : (x7 & ~x8)))) | (x4 & ~x7 & (x6 ? x5 : x8)))) | (~x3 & ((x4 & ((x5 & ~x8 & (x7 | (x6 & ~x7))) | (x7 & x8 & ~x5 & x6))) | (x7 & x8 & x5 & ~x6))) | (~x7 & ~x8 & x5 & ~x6))) | (~x4 & ((~x7 & (x3 ? (x8 & (x5 ^ ~x6)) : (x5 & ~x8))) | (x6 & x7 & x8 & ~x3 & x5))) | (~x3 & x4 & ~x5 & ~x6 & ~x8))))) | (x0 & (x7 ? ((x6 & ((x1 & ((x3 & x5 & x8) | (~x5 & ~x8 & ~x3 & x4))) | (~x5 & ((~x1 & x3 & x4 & x8) | (~x3 & ~x4 & ~x8))))) | (x1 & ~x4 & ~x6 & (x3 ? ~x8 : (x5 & x8)))) : ((~x1 & ~x3 & x6 & (x8 ? ~x5 : ~x4)) | (x1 & x3 & x4 & x5 & ~x8)))) | (~x0 & x1 & ((~x8 & (x3 ? ((~x6 & x7 & ~x4 & x5) | (x4 & ~x5 & x6 & ~x7)) : (~x5 & (x4 ? (~x6 & x7) : x6)))) | (x5 & x8 & (x3 ? (x4 & x7) : (~x4 & ~x7)))));
  assign z03 = (x2 & ((x6 & ((x7 & (x1 ? (x5 ? ((~x0 & x4 & (~x3 ^ x8)) | (x0 & ~x3 & ~x4 & x8)) : ((x4 & (x0 ? (~x8 | (x3 & x8)) : (x3 & ~x8))) | (~x0 & x3 & ~x4))) : (x0 ? (x5 & ((~x4 & ~x8) | (x3 & (x4 ^ x8)))) : (~x3 & (x4 ? (~x5 & x8) : (x5 & ~x8)))))) | (~x7 & ((x4 & (x0 ? (~x1 & (x3 ? ~x5 : (x5 & x8))) : (x3 & (x5 ^ x8)))) | (x1 & ~x3 & ((~x8 & (x0 ? (~x4 & ~x5) : (~x5 | (~x4 & x5)))) | (~x4 & x5 & x8))))) | (x1 & ((~x0 & ~x3 & x4 & x5 & x8) | (~x4 & ~x8 & x0 & x3))))) | (~x6 & (x1 ? (x3 ? (x0 ? ((x7 & x8 & x4 & x5) | (~x7 & ~x8 & ~x4 & ~x5)) : (x5 ? (x4 ? (x7 & ~x8) : ~x7) : (~x7 & ~x8))) : ((~x0 & ((~x4 & ~x7 & ~x8) | (x8 & ((x4 & (~x5 ^ x7)) | (~x5 & x7))))) | (~x4 & x7 & (x5 ^ x8)))) : ((x0 & ((~x7 & ((~x4 & x5 & ~x8) | (~x3 & (x5 | (x4 & ~x5 & ~x8))))) | (x3 & ~x4 & ~x5 & x7 & ~x8))) | (x3 & (x5 ? (x7 & x8) : ((~x4 & ~x7 & x8) | (x7 & ~x8 & ~x0 & x4))))))) | (~x0 & x1 & x3 & ~x7 & x8 & x4 & x5) | (x0 & ~x1 & ~x3 & x7 & ~x8 & ~x4 & ~x5))) | (~x2 & ((x1 & ((x0 & (x4 ? (x5 ? ((x6 & ~x7 & x8) | (x3 & x7 & ~x8)) : ((x6 & x7 & x8) | (~x7 & (x3 ? (~x6 | (x6 & ~x8)) : (~x6 & x8))))) : ((~x3 & x6 & x7 & (~x5 | (x5 & ~x8))) | (~x7 & ~x8 & x3 & x5)))) | (~x0 & (x3 ? (x4 ? (x7 & (~x8 | (x5 & ~x6 & x8))) : (x5 ? (~x7 & (x6 ^ ~x8)) : (~x6 & x8))) : (x7 & ((~x4 & x8 & (~x5 | (x5 & x6))) | (~x5 & x6 & ~x8))))) | (~x6 & ~x7 & ~x8 & ~x3 & x4 & x5))) | (x0 & ((~x3 & (x4 ? ((~x1 & ~x8 & (x5 ? (x6 & ~x7) : x7)) | (x7 & x8 & x5 & x6)) : (~x6 & ((~x5 & ~x7 & ~x8) | (~x1 & (~x7 ^ x8)))))) | (~x1 & ((x3 & ((x4 & ((x7 & x8 & ~x5 & x6) | (~x7 & ~x8 & x5 & ~x6))) | (x6 & ((x5 & x7 & x8) | (~x4 & ~x8 & (~x5 ^ ~x7)))) | (~x6 & ~x7 & ~x8 & ~x4 & ~x5))) | (x4 & ~x5 & ~x6 & ~x7 & x8))))))) | (~x3 & ((x4 & ~x7 & ((x0 & x8 & (x1 ? x6 : (x5 & ~x6))) | (~x0 & x1 & x5 & ~x6 & ~x8))) | (x0 & ~x1 & ~x4 & x7 & ~x8 & x5 & x6))) | (x3 & x8 & ((~x4 & ((x0 & ~x5 & x6 & (~x1 ^ x7)) | (~x0 & x1 & x5 & ~x6 & x7))) | (~x0 & x1 & x4 & ~x5 & ~x6 & ~x7)));
  assign z04 = (x2 & ((~x5 & (x0 ? (x7 ? ((x3 & (x1 ? (x4 ? (x6 & x8) : ~x8) : (~x4 & (x8 | (x6 & ~x8))))) | (x4 & x6 & (x1 ? ~x8 : (~x3 & x8))) | (~x4 & ~x6 & x8)) : ((x3 & ((~x4 & ~x6 & x8) | (x6 & ~x8 & ~x1 & x4))) | (~x1 & ~x3 & (x4 ? (~x6 & ~x8) : x6)))) : ((~x1 & x4 & ((~x7 & x8 & x3 & ~x6) | (x7 & ~x8 & ~x3 & x6))) | (x1 & ((x6 & ((x3 & (~x7 ^ ~x8)) | (~x4 & ((x7 & x8) | (~x3 & ~x7 & ~x8))))) | (~x3 & ~x6 & (x7 ? x8 : (~x8 | (~x4 & x8)))))) | (~x6 & ~x7 & ~x8 & x3 & ~x4)))) | (x5 & ((x1 & ((~x3 & ((x6 & ((~x0 & ((~x7 & x8) | (x4 & x7 & ~x8))) | (~x4 & ((~x7 & ~x8) | (x0 & x7 & x8))))) | (~x7 & ((x4 & ~x6 & x8) | (x0 & (x4 ? ~x8 : (~x6 & x8))))))) | (x0 & ((x4 & ~x6 & x7 & (~x8 | (x3 & x8))) | (x3 & ~x4 & x6 & (~x8 | (~x7 & x8))))) | (x4 & ~x7 & ~x8 & ~x0 & x3))) | (~x1 & ((x3 & ((x7 & (x0 ? (x4 ? (~x6 & ~x8) : (x6 & x8)) : (x4 & (~x6 | (x6 & ~x8))))) | (x0 & ~x7 & x8 & (x6 | (~x4 & ~x6))))) | (x0 & ((x6 & ((~x3 & (x4 ^ x7)) | (~x4 & x7 & ~x8))) | (~x3 & ~x6 & ~x7))) | (~x0 & ~x3 & ~x4 & x6 & x8))) | (~x3 & x4 & ~x6 & ~x7 & ~x8))) | (~x0 & x7 & ((x1 & (x3 ? (x6 & x8) : (~x4 & ~x6))) | (~x6 & ~x8 & x3 & ~x4))))) | (~x2 & ((x1 & ((x5 & ((x3 & (x0 ? (~x8 & (x6 ? (x4 | (~x4 & ~x7)) : ~x7)) : ((~x7 & x8 & ~x4 & x6) | (x4 & ~x6 & x7)))) | (~x3 & (x4 ? ((~x6 & ~x7 & ~x8) | (x7 & x8 & x0 & x6)) : (x0 ? ((~x7 & x8) | (~x6 & x7 & ~x8)) : (x6 & (~x7 ^ x8))))) | (x0 & x8 & (x4 ? (x6 & ~x7) : (~x6 & x7))))) | (x3 & ((~x5 & ((~x8 & ((x0 & x7 & (x4 | (~x4 & x6))) | (~x0 & (x4 ? x6 : (~x6 & ~x7))) | (x4 & ~x6 & ~x7))) | (x7 & x8 & ~x0 & ~x4))) | (~x0 & x4 & ~x6 & ~x7 & x8))) | (~x5 & ((~x3 & ((x8 & ((x0 & x7 & (x4 | (~x4 & x6))) | (x6 & ~x7 & (~x4 | (~x0 & x4))))) | (x7 & ~x8 & ~x0 & ~x4))) | (~x6 & x7 & ~x8 & x0 & x4))))) | (x0 & ((~x1 & ((x3 & (x8 ? ((x5 & ~x6 & x7) | (~x4 & ~x5 & x6 & ~x7)) : (x4 ? (x5 | (~x5 & x6 & x7)) : (x5 ? (x6 & x7) : (~x6 & ~x7))))) | (x4 & ~x5 & ~x6 & ~x7 & x8) | (~x3 & (x4 ? ((x6 & x7 & x8) | (x5 & ~x6 & ~x8)) : (x5 ? (x8 & (x6 ^ x7)) : (~x6 & (~x7 | ~x8))))))) | (~x3 & ((~x4 & ~x6 & ~x7 & (x5 ^ ~x8)) | (x6 & x7 & ~x8 & x4 & x5))))))) | (x0 & ~x5 & ((x8 & ((x6 & ((x1 & x3 & (x4 ^ x7)) | (~x4 & ~x7 & ~x1 & ~x3))) | (~x1 & ~x3 & ~x4 & ~x6 & x7))) | (x6 & ~x7 & ~x8 & x1 & ~x3 & x4)));
  assign z05 = (~x8 & ((x4 & (((~x5 ^ x7) & ((~x3 & x6 & x0 & ~x2) | (~x0 & ~x1 & x2 & x3 & ~x6))) | (x5 & ((x2 & ((~x0 & ((x1 & ~x3 & x7) | (x3 & x6 & ~x7))) | (~x1 & ((x0 & (x3 ? (x6 & ~x7) : (~x6 & x7))) | (x3 & x6 & x7))) | (x0 & x1 & x3 & ~x6 & ~x7))) | (x1 & ((~x2 & ((~x3 & ~x6 & ~x7) | (x0 & x3 & (x6 | (~x6 & x7))))) | (~x0 & ~x6 & (~x3 ^ x7)))) | (x0 & ~x1 & ~x2 & ~x7 & (~x3 ^ ~x6)))) | (x1 & ((~x2 & ((~x0 & x3 & (x6 ? ~x5 : ~x7)) | (~x6 & x7 & x0 & ~x5))) | (x0 & x2 & ~x5 & x7 & (x6 | (x3 & ~x6))))) | (x2 & ~x5 & x6 & (x0 ? (~x1 & ~x3) : (x3 & x7))))) | (~x4 & (x1 ? (x2 ? (x3 ? ((x6 & x7 & ~x0 & x5) | (~x6 & ~x7 & x0 & ~x5)) : ((~x6 & x7) | (~x0 & ~x7 & (x5 ^ ~x6)))) : (x0 ? (x3 ? (x5 ? (~x6 & ~x7) : (x6 & x7)) : (x5 ? (~x6 & x7) : (x6 & ~x7))) : (x3 ? (~x5 & x7) : (x5 ? ~x7 : (x6 & x7))))) : (((~x3 | (x3 & ~x7)) & ((x5 & x6 & ~x0 & x2) | (~x5 & ~x6 & x0 & ~x2))) | (x0 & ((x3 & ((x6 & ~x7) | (~x6 & x7 & x2 & x5))) | (~x3 & ((x5 & x6 & x7) | (~x2 & ~x6 & ~x7))) | (x2 & (x5 ? (~x6 ^ x7) : (~x6 & x7)))))))) | (x1 & ~x2 & ((~x0 & ~x5 & (x3 ? (~x6 & x7) : (x6 & ~x7))) | (x0 & ~x3 & x5 & x6 & ~x7))))) | (x8 & ((x2 & ((x7 & ((x0 & ((x1 & ((x3 & x4 & ~x5 & x6) | (~x3 & x5 & ~x6))) | (x3 & ((~x1 & (~x6 | (~x4 & x5 & x6))) | (~x4 & x5 & ~x6))) | (~x1 & ~x3 & x4 & ~x5 & x6))) | (~x1 & ((x4 & x6 & ~x0 & ~x3) | (x3 & ~x4 & x5 & ~x6))) | (~x0 & ((x1 & ~x4 & (~x3 ^ x6)) | (x5 & x6 & x3 & x4))) | (x1 & ~x3 & x4 & ~x5 & ~x6))) | (~x0 & ((x4 & ((x1 & (x3 ? (~x5 & ~x7) : (x5 & x6))) | (~x1 & ~x3 & ~x5 & x6 & ~x7))) | (~x1 & x3 & x5 & ~x6 & ~x7))) | (~x7 & ((x0 & ((~x3 & ((x1 & x5 & (x4 ^ x6)) | (~x5 & x6 & ~x1 & ~x4))) | (~x4 & ((~x1 & x5 & x6) | (x3 & ~x5 & ~x6))))) | (~x1 & x3 & ~x4 & ~x5 & ~x6))))) | (~x2 & ((x1 & (x0 ? ((~x7 & ((x4 & ((x5 & x6) | (~x3 & ~x5 & ~x6))) | (x3 & x5 & ~x6))) | (~x5 & ((x3 & (x4 ? (~x6 & x7) : x6)) | (x4 & x6 & x7)))) : ((x3 & ((x4 & ~x7) | (~x6 & x7 & ~x4 & ~x5))) | (x7 & ((~x3 & (x4 ? (~x5 & x6) : x5)) | (x4 & x5 & x6))) | (~x6 & ~x7 & ~x3 & ~x5)))) | (x0 & ((x5 & ((x3 & ((x4 & ~x6 & x7) | (x6 & ~x7 & ~x1 & ~x4))) | (~x1 & x7 & ((~x4 & x6) | (x4 & ~x6) | (~x3 & (x4 ^ ~x6)))))) | (~x1 & x4 & ((x6 & ~x7) | (~x6 & x7 & ~x3 & ~x5))) | (~x3 & ~x4 & ~x5 & x6 & x7))))) | (x0 & ~x6 & ((~x1 & ~x3 & (x4 ? (x5 & ~x7) : (~x5 & x7))) | (x1 & x3 & ~x4 & ~x5 & x7))))) | (x0 & ((x2 & ((x6 & ((x3 & ((~x4 & x5 & ~x7) | (x1 & ~x5 & (x4 ^ x7)))) | (~x1 & ~x3 & ~x4 & x5 & x7))) | (~x1 & ~x3 & x5 & ~x6 & ~x7))) | (x1 & ~x2 & x3 & ~x6 & ~x7 & x4 & ~x5))) | (~x0 & x1 & x3 & x6 & ((~x2 & (x4 ? (~x5 & x7) : x5)) | (~x5 & ~x7 & x2 & ~x4)));
  assign z06 = (x2 & ((~x8 & (x1 ? (x0 ? (x3 ? ((x4 & (x6 ? ~x5 : x7)) | (x5 & x6 & ~x7) | (~x4 & (x6 | (~x5 & (x7 | (~x6 & ~x7)))))) : ((x4 & x6 & x7) | (~x6 & ~x7 & ~x4 & x5))) : (x6 ? ((~x4 & ~x5 & ~x7) | (x3 & x7 & (x5 | (x4 & ~x5)))) : (x3 ? (x5 & ~x7) : (x4 ? x7 : (~x5 & ~x7))))) : ((~x7 & ((x3 & ((~x4 & x5 & x6) | (~x0 & (x4 ? x5 : (~x5 & ~x6))))) | (~x3 & ((x0 & ~x6 & (x5 | (x4 & ~x5))) | (~x5 & x6 & ~x0 & x4))) | (x0 & ~x5 & x6))) | (~x0 & ((x3 & ~x4 & x5 & ~x6) | (x4 & x6 & x7))) | (x0 & ((~x4 & ~x5 & ~x6) | (x7 & ((x3 & (x4 ? (x5 & ~x6) : (~x5 & x6))) | (x6 & (~x3 | (~x4 & x5)))))))))) | (x8 & ((x6 & ((x1 & ((x3 & ((x0 & ~x5 & (~x4 ^ x7)) | (~x4 & x5 & ~x7) | (~x0 & x4 & x7))) | (~x0 & ~x3 & x5 & (x4 | x7)))) | (~x1 & ((~x3 & ((x0 & ~x5 & (~x4 | (x4 & x7))) | (x5 & ~x7 & ~x0 & ~x4))) | (x5 & x7 & ~x0 & x3))) | (~x0 & x3 & x4 & ~x5 & ~x7))) | (~x6 & (x0 ? (~x7 & ((~x3 & x4 & x5) | (~x4 & (x5 ? x1 : x3)))) : ((x4 & ((x3 & (x1 ? (~x5 & ~x7) : (x7 | (x5 & ~x7)))) | (x1 & ((~x5 & x7) | (~x3 & x5 & ~x7))))) | (~x3 & ~x4 & x5 & x7)))) | (~x4 & x5 & ~x7 & ~x0 & x1 & ~x3))) | (x5 & ((x3 & x4 & ((x0 & (x1 ? (x6 & x7) : (~x6 & ~x7))) | (x6 & ~x7 & ~x0 & x1))) | (x0 & ~x1 & ~x3 & ~x4 & x6 & x7))) | (~x0 & x1 & ~x4 & x7 & (x3 ? (~x5 & x6) : ~x6)))) | (x1 & ((~x0 & ((~x3 & (x4 ? ((~x7 & ~x8 & x5 & ~x6) | (x6 & x7 & ~x2 & ~x5)) : ((x6 & (x5 ? (~x7 & ~x8) : (x7 & (~x8 | (~x2 & x8))))) | (~x2 & x5 & ~x6 & (~x8 | (x7 & x8)))))) | (~x2 & ((x3 & ((~x4 & (x5 ? ~x7 : (~x6 & x8))) | (~x8 & ((~x5 & (x6 ? x4 : x7)) | (x4 & (~x6 ^ x7)))) | (~x7 & x8 & (x5 ? x4 : x6)))) | (x6 & x7 & x8 & ~x4 & x5))))) | (x0 & ((~x2 & ((x3 & ((~x4 & x6 & (x5 ? x8 : x7)) | (~x6 & ((x5 & ~x8 & (~x7 | (x4 & x7))) | (x4 & ~x5 & (~x7 | (x7 & x8))))))) | (x4 & ((x5 & x6 & (x7 ? ~x3 : x8)) | (~x3 & x7 & (x8 ? ~x5 : ~x6)))) | (~x6 & x7 & ~x8 & ~x3 & ~x4 & x5))) | (~x3 & ((x4 & ~x5 & (x7 ? ~x8 : x6)) | (x7 & x8 & ~x4 & x6))) | (x6 & ~x7 & x8 & x3 & x4 & ~x5))) | (x8 & ((~x6 & x7 & ~x4 & ~x5) | (~x2 & ((~x3 & ~x5 & ~x7 & (x4 ^ x6)) | (x3 & x5 & ~x6 & x7))))))) | (x0 & ((~x4 & (x8 ? ((~x5 & ((~x1 & ~x3 & x7 & (~x6 | (~x2 & x6))) | (x6 & ~x7 & ~x2 & x3))) | (~x1 & x5 & ~x6 & (x7 | (x3 & ~x7)))) : ((~x1 & ((x5 & x7 & (x6 ? ~x3 : ~x2)) | (~x2 & ~x3 & ~x6 & (~x5 | ~x7)))) | (~x2 & ~x3 & ~x5 & (~x6 ^ x7))))) | (~x1 & ((~x2 & ((x4 & (x3 ? ((~x7 & ~x8 & x5 & ~x6) | (~x5 & (x6 ? (~x8 | (x7 & x8)) : (~x7 & x8)))) : (x5 ? (x7 & (x6 ^ ~x8)) : (x6 & x8)))) | (x6 & ~x7 & x8 & ~x3 & x5))) | (x6 & ~x7 & ~x8 & ~x3 & x4 & x5))) | (x7 & x8 & x5 & ~x6 & ~x2 & x3 & x4)));
  assign z07 = (~x8 & (x0 ? ((x5 & (x1 ? ((~x3 & ((x6 & x7 & ~x2 & ~x4) | (x2 & ~x7))) | (x2 & ((x4 & ~x6 & x7) | (x3 & x6 & ~x7)))) : (x4 ? (x3 ? (x7 ? ~x2 : x6) : ((~x6 & x7) | (x2 & x6 & ~x7))) : ((~x6 & (x2 ? (~x7 | (x3 & x7)) : x7)) | (~x2 & x3 & x6))))) | (~x5 & (x2 ? ((x3 & (x7 ? ((x4 & ~x6) | (~x1 & ~x4 & x6)) : ((~x4 & x6) | (x1 & (x4 ^ ~x6))))) | (~x1 & ~x3 & ((~x6 & x7) | (x4 & (x6 | (~x6 & ~x7)))))) : ((x1 & x4 & (x3 ? ~x7 : x6)) | (~x3 & ~x4 & (x6 ? x7 : (~x1 | ~x7)))))) | (x2 & ((x1 & x3 & (x4 ? (~x6 & ~x7) : x6)) | (x6 & x7 & ~x1 & ~x3))) | (~x4 & ~x6 & ~x7 & ~x1 & ~x2 & ~x3)) : ((x3 & ((x2 & ((x5 & ((~x1 & (x7 ? x6 : x4)) | (x4 & (x6 ? x1 : x7)))) | (x6 & x7 & x4 & ~x5))) | (x1 & ~x2 & ((~x5 & (~x4 | (x4 & x6))) | (x4 & ~x6 & (x7 | (x5 & ~x7))))))) | (x1 & ((~x6 & x7 & ~x4 & ~x5) | (~x3 & ((x2 & (x4 ? (~x5 & x7) : (~x6 & ~x7))) | (x4 & ((x5 & ~x6 & ~x7) | (~x2 & x6 & x7))) | (~x4 & ((~x5 & x6) | (~x2 & x5 & (~x6 | (x6 & ~x7))))))))) | (x5 & x6 & ~x7 & ~x1 & x2 & ~x4)))) | (x8 & ((x6 & ((x4 & ((x0 & ((~x2 & (x1 ? ((~x5 & (x7 | (x3 & ~x7))) | (~x3 & x5 & x7)) : (x3 ? x7 : (~x5 & ~x7)))) | (x1 & ~x3 & ~x7))) | (~x0 & ((x5 & (x1 ? (x2 ^ x3) : (x2 & x7))) | (x2 & ~x7 & (x3 ? ~x5 : ~x1)))) | (x3 & ~x5 & x7 & x1 & x2))) | (~x4 & ((x0 & (x1 ? ((x5 & x7 & x2 & ~x3) | (~x2 & x3 & ~x7)) : ((~x3 & ~x5) | (~x2 & x5 & ~x7)))) | (~x0 & ((x2 & ((x3 & ~x5 & x7) | (x1 & ~x3 & x5 & ~x7))) | (x1 & ~x2 & ((~x5 & x7) | (x3 & x5 & ~x7))))) | (x3 & ~x5 & ~x7 & x1 & x2))) | (~x3 & x5 & x7 & ~x0 & x1 & x2))) | (~x6 & ((x2 & ((~x0 & ((x1 & x4 & ~x5) | (~x3 & ~x4 & x5 & ~x7))) | (~x1 & x3 & x5 & (~x4 ^ x7)) | (~x4 & ~x5 & ~x7 & x0 & x1 & ~x3))) | (~x2 & ((x1 & ((x3 & ((~x5 & (x0 ? (~x4 ^ x7) : ~x4)) | (~x0 & x5 & ~x7))) | (x0 & ((~x4 & x5 & x7) | (~x3 & x4 & ~x5 & ~x7))))) | (x0 & ~x1 & (x3 ? (~x5 & (x4 ^ x7)) : (x4 & x7))))) | (x0 & ((x1 & x3 & ~x4 & ~x5 & x7) | (~x1 & ~x3 & x4 & x5 & ~x7))))) | (x1 & ~x2 & ((~x0 & ((~x4 & x5 & x7) | (~x3 & x4 & ~x5))) | (~x4 & x5 & ~x7 & x0 & ~x3))) | (x0 & ~x1 & x2 & x3 & ~x7 & (~x4 ^ x5)))) | (x0 & ~x2 & ((~x1 & ~x3 & x4 & ~x5 & x6 & x7) | (x1 & x3 & x5 & ~x6 & ~x7))) | (x2 & ~x6 & x7 & ((~x0 & ((~x3 & ~x4 & x5) | (~x1 & x4 & ~x5))) | (x1 & ~x3 & ~x4 & x5)));
  assign z08 = (x2 & ((x8 & ((~x0 & (x5 ? ((~x6 & x7 & ~x1 & x4) | (~x4 & ~x7 & x1 & ~x3)) : (x1 ? (x6 & ((~x4 & x7) | (~x3 & x4 & ~x7))) : (x3 ? (x4 & ~x7) : (x4 ? ~x6 : x7))))) | (x3 & ((~x5 & ((x6 & ((x0 & ~x7 & (~x4 | (x1 & x4))) | (x1 & x4 & x7))) | (~x4 & x7 & x0 & ~x1))) | (~x6 & ~x7 & ((x0 & ~x4) | (~x1 & x4 & x5))))) | (x0 & ((~x5 & ((~x1 & x6 & x7 & (x4 | (~x3 & ~x4))) | (x1 & ~x3 & ~x4 & ~x6 & ~x7))) | (~x3 & x5 & ((~x4 & ~x6 & x7) | (x1 & (x4 ? (~x6 & ~x7) : x6)))))) | (x1 & ~x3 & x4 & ~x5 & ~x6 & x7))) | (~x8 & ((x4 & ((~x0 & ((x6 & (x1 ? (x3 ? (~x5 & x7) : ~x7) : (x5 & x7))) | (x3 & x5 & ~x6 & x7) | (~x5 & ~x7 & ~x1 & ~x3))) | (~x7 & ((x5 & x6 & ~x1 & ~x3) | (x0 & x1 & x3 & ~x5 & ~x6))) | (x0 & ((x7 & ((x1 & (x6 ? ~x3 : x5)) | (x5 & x6 & ~x1 & x3))) | (~x5 & ~x6 & ~x1 & ~x3))) | (~x1 & x3 & ~x5 & ~x6 & x7))) | (~x7 & (x1 ? (~x3 & ((~x4 & x5 & ~x6) | (~x0 & ~x5 & (~x6 | (~x4 & x6))))) : ((x0 & (x3 ? (x5 & x6) : (~x4 & ~x5))) | (~x4 & x5 & (~x6 | (~x0 & x3 & x6)))))) | (~x4 & ((x7 & (x0 ? (x1 ? (~x5 & (x3 | (~x3 & x6))) : (x3 & ~x6)) : (x3 ? (~x5 & x6) : (x5 & ~x6)))) | (x0 & x1 & x3 & x5 & x6))))) | (~x0 & x6 & ((~x1 & ~x3 & ~x4) | (x5 & ~x7 & x1 & x3))))) | (~x2 & ((x5 & (x0 ? (x1 ? ((~x6 & ((x3 & (x8 ? x4 : ~x7)) | (~x4 & x7 & x8))) | (~x3 & x7 & (x4 ? (x6 & x8) : ~x8))) : (((x6 ? (~x7 & x8) : ~x8) & (x3 ^ x4)) | (x3 & ((x6 & x7 & x8) | (x4 & ~x7 & ~x8))) | (x7 & x8 & x4 & ~x6))) : (x1 & ((x3 & (x4 ? (x6 ? (x7 & x8) : (~x7 & ~x8)) : (~x7 & x8))) | (x6 & ((~x4 & x7 & x8) | (~x3 & ~x8 & (x7 | (~x4 & ~x7))))) | (~x3 & ~x6 & (x7 | (x4 & ~x7))))))) | (~x5 & (x0 ? ((x3 & ((x8 & ((~x1 & (x4 ? ~x7 : (~x6 & x7))) | (~x6 & ~x7 & x1 & ~x4))) | (x1 & ((x4 & ~x6 & ~x7) | (~x8 & (x4 ? (x7 | (x6 & ~x7)) : (x6 & x7))))))) | (~x3 & ((x1 & ((x4 & x7 & x8) | (~x7 & ~x8 & ~x4 & x6))) | (~x6 & ((~x4 & ~x7 & ~x8) | (~x1 & (x4 ? (x7 & x8) : ~x8)))) | (x7 & ~x8 & x4 & x6))) | (x6 & x7 & x8 & x1 & x4)) : (x1 & ((x8 & ((~x4 & (x7 | (~x3 & x6 & ~x7))) | (x3 & x6 & ~x7) | (~x3 & ~x6 & (~x7 | (x4 & x7))))) | (x6 & x7 & ~x8 & ~x3 & ~x4))))) | (x7 & ((x0 & ~x3 & ((~x4 & x6 & x8) | (~x6 & ~x8 & x1 & x4))) | (~x0 & x1 & x3 & x4 & ~x8))) | (~x0 & x1 & x3 & ~x7 & ~x8 & ~x4 & x6))) | (x4 & ~x7 & ((x1 & ((~x0 & ~x6 & ~x8 & (~x3 ^ ~x5)) | (x6 & x8 & ~x3 & x5))) | (x0 & ~x1 & ~x3 & x5 & ~x6 & x8))) | (x0 & ~x1 & ~x3 & ~x4 & x7 & (x5 ? (x6 & ~x8) : (~x6 & x8)));
  assign z09 = (~x5 & ((~x4 & (x3 ? (((x6 ? ~x8 : x7) & (x0 ? (~x1 & ~x2) : (x1 & x2))) | (x0 & ((x1 & ((~x2 & (x7 ? x6 : x8)) | (x7 & x8 & x2 & ~x6))) | (x2 & (x7 ? ~x8 : ((x6 & ~x8) | (~x1 & ~x6 & x8)))))) | (~x0 & ((x1 & ((~x6 & ~x7 & ~x8) | (~x2 & (x6 ? ~x7 : x8)))) | (x7 & x8 & x2 & x6)))) : ((x1 & ((x2 & ((~x6 & ~x8) | (x0 & x6 & x7))) | (~x8 & ((x0 & ((x6 & ~x7) | (~x2 & ~x6 & x7))) | (x6 & ~x7 & ~x0 & ~x2))) | (~x0 & x6 & x8 & (~x7 | (~x2 & x7))))) | (~x1 & ((x2 & (x0 ? (x6 & ~x7) : (x6 | (x7 & x8)))) | (x0 & ((x6 & ~x7 & x8) | (~x2 & (x6 ? (x7 & x8) : ~x8)))))) | (x0 & ~x2 & ~x8 & (~x6 ^ x7))))) | (x4 & ((x1 & ((~x0 & ((~x3 & (x8 ? ~x2 : ((x6 & ~x7) | (x2 & ~x6 & x7)))) | (x3 & ((x7 & x8 & x2 & x6) | (~x2 & (x6 ? x7 : (~x7 & x8))))) | (x2 & x8 & (x6 ^ x7)))) | (x0 & ((x6 & (x2 ? (x3 & x7) : (~x3 & ~x7))) | (~x7 & (x2 ? (~x3 ^ ~x8) : (x3 & ~x6))) | (x7 & x8 & ~x2 & ~x3))) | (~x6 & x7 & (x2 ? (~x3 & x8) : x3)))) | (x2 & ((~x1 & ((x0 & ((x6 & x7 & x8) | (~x7 & ~x8 & ~x3 & ~x6))) | (~x6 & ~x7 & ~x0 & x3))) | (x6 & x7 & x8 & ~x0 & ~x3))) | (x0 & ((~x1 & ((x8 & ((x3 & ~x6) | (~x2 & x6 & (~x3 | (x3 & x7))))) | (x7 & ~x8 & ~x3 & ~x6))) | (~x7 & x8 & x3 & x6))))) | (x6 & ((~x0 & ((~x7 & x8 & ~x1 & x2) | (x1 & ~x2 & ~x3 & x7 & ~x8))) | (~x1 & x2 & ~x3 & x7 & ~x8))))) | (x2 & ((~x6 & ((~x0 & ((x8 & ((x1 & (x3 ? (x5 & x7) : (x4 & ~x7))) | (~x1 & x3 & x4 & x5 & ~x7))) | (x5 & ((~x1 & (x3 ? (x4 & ~x8) : (~x7 & (x4 | (~x4 & ~x8))))) | (x7 & ~x8 & ~x3 & ~x4))))) | (x0 & ((~x7 & ((~x3 & (x1 ? (~x4 & (x8 | (x5 & ~x8))) : (x5 & (~x8 | (x4 & x8))))) | (x4 & x5 & ~x1 & x3))) | (x3 & ((~x8 & (x1 ? (x4 & x5) : (x7 & (x4 | (~x4 & x5))))) | (~x1 & x7 & x8))))) | (~x3 & x5 & x7 & (x1 ? ~x4 : (x4 & ~x8))))) | (x6 & ((x1 & ((~x4 & (x0 ? ((x3 & ~x8) | (x7 & x8 & ~x3 & x5)) : (x7 & (x3 ? x8 : (x5 & ~x8))))) | (~x0 & x4 & x5 & (x3 ? ~x7 : x8)))) | (~x0 & ((~x1 & ~x7 & ((~x3 & x4) | (x3 & ~x4 & x5 & ~x8))) | (x7 & ~x8 & x3 & x4))) | (x5 & ~x7 & ~x8 & x0 & ~x1 & x4))) | (~x4 & x5 & ~x7 & ~x0 & x1 & x3))) | (x5 & ((~x2 & ((x3 & (x0 ? ((~x8 & ((~x4 & (x1 ? (~x6 & ~x7) : (~x6 | (x6 & ~x7)))) | (x1 & x4 & (x6 ^ x7)))) | (~x6 & x8 & (~x4 | (x1 & ~x7)))) : (x1 & ((~x4 & ~x7 & x8) | (~x6 & (x4 ? (~x7 ^ x8) : ~x8)))))) | (x7 & (x0 ? (~x1 & ~x6 & ((~x4 & ~x8) | (~x3 & x4 & x8))) : (x1 & ~x3 & (x4 ? x6 : x8)))) | (~x8 & ((~x0 & x1 & ~x7 & (x4 ? x6 : ~x3)) | (x0 & ~x1 & ~x3 & x4 & x6))))) | (x0 & ~x1 & ~x4 & x6 & (x3 ? (~x7 & x8) : (x7 & ~x8))) | (~x0 & x1 & ~x3 & ~x7 & ~x8 & x4 & ~x6))) | (x0 & ~x2 & ~x3 & x8 & ((x1 & x4 & x6) | (~x6 & x7 & ~x1 & ~x4)));
  assign z10 = (x3 & ((~x2 & (((x8 | (~x6 & ~x8)) & ((~x4 & ~x5 & x7 & x0 & ~x1) | (~x0 & x1 & x4 & x5 & ~x7))) | (x0 & ((~x1 & ((x8 & ((x4 & ((~x6 & ~x7) | (~x5 & x6 & x7))) | (x5 & ((~x6 & x7) | (~x4 & x6 & ~x7))))) | (x6 & ~x7 & ~x8 & ~x4 & ~x5))) | (~x8 & ((x4 & ~x6 & ((~x5 & ~x7) | (x1 & x5 & x7))) | (x1 & ~x4 & (x5 ? x7 : (~x7 | (x6 & x7)))))) | (~x6 & ~x7 & x8 & x1 & x5))) | (~x5 & x7 & ~x8 & ~x0 & x1 & ~x4))) | (x2 & ((x1 & (x6 ? (x0 ? ((~x4 & (x5 ^ x8)) | (~x7 & x8 & (x5 | (x4 & ~x5)))) : (x4 & (x5 ? (~x7 | (x7 & x8)) : (x7 & ~x8)))) : ((~x0 & ((x4 & ~x5 & x7) | (x5 & ~x7 & ~x8))) | (x0 & x5 & ~x7) | (x7 & x8 & x4 & ~x5)))) | (~x1 & (x5 ? (x8 ? ((x4 & ~x6 & ~x7) | (~x0 & x6 & x7)) : (x0 ? ((~x6 & x7) | (x4 & x6 & ~x7)) : (~x7 & (x4 ^ x6)))) : ((~x0 & ~x4 & (x7 ? ~x6 : ~x8)) | (x7 & ~x8 & x0 & x4)))) | (~x5 & ((~x0 & ~x8 & (x4 ? (~x6 & ~x7) : (x6 & x7))) | (~x7 & x8 & ~x4 & ~x6))) | (~x6 & x7 & x8 & x0 & ~x4 & x5))) | (x0 & ~x6 & ((~x5 & x8 & ~x1 & x4) | (x7 & ~x8 & x1 & ~x4))) | (~x0 & x1 & ~x5 & x6 & ~x7 & (x4 ^ x8)))) | (~x3 & ((x0 & ((x6 & ((~x8 & ((~x1 & ~x7 & (~x4 | (~x2 & x4 & x5))) | (x1 & ((~x2 & x4 & (x5 | (~x5 & x7))) | (x5 & x7 & x2 & ~x4))) | (~x5 & x7 & ~x2 & ~x4))) | (x8 & ((x7 & (x1 ? (x2 ? x4 : x5) : (x2 ? (~x4 & ~x5) : (x4 & x5)))) | (x2 & ~x5 & (x1 ? ~x7 : x4)))) | (x1 & x2 & x4 & x5 & x7))) | (~x6 & ((x1 & (x2 ? (~x7 & ((x5 & x8) | (~x4 & (~x5 | (x5 & ~x8))))) : (~x8 | (x4 & x7)))) | (~x1 & ((x2 & ((x7 & x8) | (~x7 & ~x8 & x4 & ~x5))) | (~x4 & ~x5 & (~x7 | (x7 & x8))))) | (~x5 & ~x8 & ~x2 & x4))) | (~x1 & ~x4 & x5 & (x7 ? x2 : x8)))) | (x2 & ((~x6 & ((~x5 & ((x7 & ~x8 & x1 & ~x4) | (x4 & x8 & ~x0 & ~x1))) | (~x0 & ((x1 & x7 & (x4 ^ x8)) | (x5 & ~x7 & ((~x4 & x8) | (~x1 & (x4 | (~x4 & ~x8))))))) | (x5 & x7 & ~x8 & ~x1 & x4))) | (~x0 & ((x8 & ((x1 & ((x5 & x6 & x7) | (x4 & ~x5 & ~x7))) | (x6 & ~x7 & ~x1 & x4))) | (~x1 & x4 & ~x5 & x6 & (x7 | (~x7 & ~x8))))))) | (x1 & ((~x0 & ((~x2 & ((~x5 & ((x4 & (x7 ? x8 : x6)) | (x7 & ((~x6 & ~x8) | (~x4 & x6 & x8))))) | (~x4 & x5 & ((~x6 & ~x8) | (~x7 & (x8 | (x6 & ~x8))))))) | (x7 & ~x8 & ~x5 & x6))) | (~x6 & ~x7 & ~x8 & ~x2 & ~x5))))) | (x5 & ((x7 & ((x6 & ((~x0 & ((x1 & ~x2 & ~x4) | (~x1 & x2 & x4 & ~x8))) | (~x1 & x2 & ((x4 & x8) | (x0 & ~x4 & ~x8))))) | (x0 & ~x1 & ~x2 & ~x6 & (~x4 ^ x8)) | (~x4 & x8 & x1 & x2))) | (x1 & ~x7 & ((x4 & x8 & x0 & ~x2) | (~x0 & x2 & ~x4 & x6 & ~x8))))) | (x0 & x2 & x4 & ~x7 & x8 & ~x5 & ~x6);
  assign z11 = (x6 & ((x2 & (x5 ? ((~x0 & ((x4 & (x1 ? (~x3 & ~x7) : (x3 ? (x7 & x8) : (~x7 & ~x8)))) | (x3 & ~x4 & (x7 ? ~x8 : ~x1)))) | (x0 & ((x1 & x4 & x7) | (x8 & (x1 ? (x3 ? (x4 & ~x7) : (~x4 & x7)) : (x3 ? (~x4 & x7) : (x4 & ~x7)))))) | (~x7 & ~x8 & ~x3 & ~x4)) : (((~x7 ^ ~x8) & ((~x0 & ~x3 & x4) | (x3 & ~x4 & x0 & x1))) | (~x1 & (x0 ? (x3 ? (x4 & x7) : (~x4 & ~x7)) : (x4 ? (~x7 & ~x8) : ~x3)))))) | (~x2 & ((x1 & (x3 ? ((~x5 & ((~x4 & x7 & x8) | (~x0 & (x4 ? x7 : (~x7 & ~x8))))) | (~x0 & x4 & ((x7 & ~x8) | (x5 & ~x7 & x8)))) : ((x0 & ((~x4 & x5 & x7) | (~x7 & (x4 ? (~x5 | (x5 & ~x8)) : (~x5 & x8))))) | (~x0 & ~x4 & x5 & ~x7 & ~x8)))) | (x0 & ((x7 & ((~x3 & ((x4 & ~x5 & ~x8) | (~x1 & x8 & (~x4 ^ x5)))) | (~x1 & x3 & ~x4 & ~x5))) | (~x1 & x3 & ~x4 & ~x7 & (x5 | (~x5 & x8))))))) | (~x7 & ~x8 & x4 & ~x5 & x0 & x1 & x3))) | (~x6 & ((~x1 & (x0 ? ((~x7 & (x2 ? ((x4 & ~x5 & x8) | (x3 & ((~x5 & ~x8) | (~x4 & x5 & x8)))) : ((~x3 & ~x4 & ~x5) | (~x8 & (x3 ? (~x4 ^ x5) : ~x4))))) | (~x3 & ((x7 & ((x2 & (x4 ? (~x5 & ~x8) : x5)) | (~x5 & x8 & ~x2 & x4))) | (~x5 & ~x8 & ~x2 & ~x4))) | (x5 & x7 & ~x8 & x2 & x3 & ~x4)) : ((~x3 & ~x4) | (~x5 & x7 & x8 & x2 & x3 & x4)))) | (x1 & ((x7 & (x0 ? (~x2 & ((x3 & ((x5 & ~x8) | (x4 & ~x5 & x8))) | (x4 & x5 & x8) | (~x5 & ~x8 & ~x3 & ~x4))) : (x2 ? (x3 & (~x4 ^ x5)) : (~x3 & ((~x4 & x5 & x8) | (~x5 & (~x8 | (x4 & x8)))))))) | (~x7 & ((x4 & ((x2 & ((x0 & ~x3 & x5) | (x3 & ~x5 & x8))) | (~x0 & ~x2 & ((~x3 & x5) | (~x5 & x8) | (x3 & ~x8))))) | (x0 & x2 & ~x4 & ~x5 & (~x8 | (~x3 & x8))))) | (x4 & x5 & x8 & x0 & ~x2 & x3))) | (x5 & x8 & ((~x0 & x2 & ~x3 & (~x4 ^ x7)) | (x3 & x4 & x7 & x0 & ~x2))))) | (~x0 & ~x1 & ~x2);
  assign z12 = (x1 & ((~x4 & ((x5 & (x8 ? ((x7 & ((x0 & (x6 ? ~x2 : ~x3)) | (~x3 & ~x6 & ~x0 & ~x2))) | (x6 & ~x7 & ~x0 & x3)) : ((~x3 & (x0 ? (x2 ? ~x7 : (x6 & x7)) : (~x6 & ~x7))) | (~x0 & (x2 ? (x3 & x7) : (x6 & ~x7)))))) | (~x2 & ((~x5 & ((x0 & ((x3 & x6 & x7) | (~x7 & x8 & ~x3 & ~x6))) | (~x0 & ((x7 & x8 & ~x3 & x6) | (x3 & ~x7 & ~x8))) | (x7 & x8 & x3 & ~x6))) | (~x6 & x7 & ~x8 & x0 & ~x3))))) | (x4 & ((x3 & ((~x5 & ((~x6 & ((x0 & (x2 ? (~x7 & ~x8) : (x7 & x8))) | (~x2 & ~x7 & (~x8 | (~x0 & x8))))) | (x6 & x7 & ~x0 & x2))) | (x2 & ((x0 & ((~x6 & ~x7 & x8) | (x5 & x6 & x7))) | (x7 & ~x8 & x5 & ~x6))))) | (x2 & ~x3 & ((~x7 & ((x0 & (x5 ^ x6)) | (~x0 & ~x5 & ~x6 & x8))) | (x7 & ~x8 & ~x0 & ~x5))))) | (x2 & x6 & ~x7 & x8 & (x0 ? (x3 & x5) : (~x3 & ~x5))))) | (~x1 & (x0 ? (x4 ? ((x5 & ((x2 & ((x7 & ~x8 & x3 & x6) | (~x3 & ~x7 & x8))) | (~x2 & ((~x3 & x7 & x8) | (~x7 & ~x8 & x3 & ~x6))) | (~x7 & ~x8 & ~x3 & x6))) | (~x2 & ~x5 & x7 & (x3 ? (x6 & x8) : ~x6))) : (x2 ? ((~x5 & ((~x7 & ((x6 & x8) | (~x3 & (~x6 | ~x8)))) | (x7 & ~x8 & x3 & x6))) | (x3 & x5 & ~x6 & (~x7 ^ ~x8))) : ((x6 & x7 & x8 & ~x3 & x5) | (~x6 & ~x7 & ~x8 & x3 & ~x5)))) : ((x2 & ((x5 & ((~x7 & ~x8 & ~x4 & x6) | (x3 & (x4 ? (x6 & x7) : (~x6 & ~x7))))) | (~x3 & ~x5 & (x4 ? (~x7 & ~x8) : x6)))) | ~x2 | (~x3 & ~x6 & (~x4 | (~x5 & ~x7 & x8)))))) | (~x0 & x2 & x5 & ~x6 & x8 & (x3 ? (x4 & x7) : (~x4 & ~x7))) | (x3 & x4 & x0 & ~x2 & ~x7 & ~x8 & ~x5 & x6);
  assign z13 = (x0 & ((~x3 & (((x4 ? (x5 & x8) : ~x5) & ((x6 & x7 & x1 & ~x2) | (~x6 & ~x7 & ~x1 & x2))) | (~x2 & ((~x1 & ((x4 & (x5 ? (~x7 & ~x8) : (x6 & x7))) | (x7 & x8 & ~x4 & x5))) | (x6 & ~x7 & x8 & x1 & ~x4 & ~x5))) | (x1 & x2 & ((~x7 & ~x8 & x4 & ~x5) | (~x4 & ((~x7 & ~x8 & ~x5 & x6) | (x5 & (x6 ? (x7 & x8) : (~x7 & ~x8))))))))) | (x2 & ((x3 & (x5 ? ((x1 & ~x7 & x8 & (~x6 | (~x4 & x6))) | (x4 & x7 & ~x8 & (~x6 | (~x1 & x6)))) : ((~x1 & ~x4 & (~x7 ^ ~x8)) | (x6 & ~x8 & x1 & x4)))) | (~x5 & ~x7 & ((x6 & x8 & x1 & x4) | (~x6 & ~x8 & ~x1 & ~x4))))) | (~x2 & ((x3 & ((x8 & ((x1 & ~x4 & x7 & (x5 ^ ~x6)) | (x5 & x6 & ~x7 & ~x1 & x4))) | (x4 & ~x7 & ~x8 & (x6 ? ~x1 : ~x5)))) | (x5 & ~x6 & x7 & (x1 ? ~x4 : (x4 & x8))))))) | (~x0 & ((x2 & ((~x1 & ((~x6 & ((x4 & ((x7 & x8 & x3 & x5) | (~x7 & ~x8 & ~x3 & ~x5))) | (~x7 & ~x8 & ~x4 & x5))) | (~x4 & x6 & ((~x3 & ~x5) | (~x7 & (x3 ? (x5 ^ ~x8) : (x5 & ~x8))))))) | (x1 & ((~x5 & (x3 ? ((x6 & x7 & ~x8) | (x4 & ~x6 & (x7 | (~x7 & x8)))) : ((~x4 & ~x7 & x8) | (x7 & ~x8 & x4 & ~x6)))) | (~x4 & x5 & ((x7 & ~x8 & x3 & ~x6) | (~x3 & x6 & (~x8 | (~x7 & x8))))))) | (x6 & x7 & x8 & x3 & x4 & ~x5))) | (~x1 & (~x2 | (~x5 & ~x6 & ~x3 & ~x4))) | (x1 & ~x2 & ((x6 & ~x7 & ~x8 & ~x3 & x4 & x5) | (~x4 & ((~x7 & ((x3 & (x5 ? x8 : (~x6 & ~x8))) | (~x8 & ((x5 & ~x6) | (~x3 & ~x5 & x6))))) | (~x5 & x7 & (x6 ? x8 : ~x3)))))))) | (~x7 & ((x1 & ((~x5 & ~x6 & x8 & x2 & ~x3 & x4) | (x5 & x6 & ~x8 & ~x2 & x3 & ~x4))) | (~x1 & x2 & ~x3 & x4 & ~x5 & x6 & x8)));
  assign z14 = (x1 & ((~x7 & ((x3 & (((x6 ^ ~x8) & ((x4 & x5 & ~x0 & ~x2) | (x0 & x2 & ~x5))) | (~x4 & x5 & ~x6 & (x0 ? (x2 & x8) : ~x2)))) | (~x3 & (x5 ? ((~x0 & (x2 ? (x4 ? x6 : (~x6 & ~x8)) : (x4 & ~x6))) | (x6 & ~x8 & ~x2 & x4)) : ((~x2 & (x0 ? (x4 & x6) : (x4 ? (~x6 & x8) : (x6 & ~x8)))) | (~x4 & ((x0 & (x8 ? ~x6 : x2)) | (~x6 & x8 & ~x0 & x2))) | (x4 & ~x6 & x0 & x2)))) | (~x0 & x2 & ~x4 & x5 & x6 & x8))) | (x7 & (x2 ? ((x6 & ((x0 & x4 & (x3 ? (~x5 & ~x8) : x5)) | (~x4 & ~x8 & ((x3 & ~x5) | (~x0 & ~x3 & x5))))) | (~x5 & ~x6 & ~x0 & x3)) : (x0 ? ((x6 & ((~x3 & (x4 ? (x5 ^ ~x8) : ~x5)) | (~x5 & ~x8 & x3 & ~x4))) | (x5 & ~x6 & ((x4 & x8) | (x3 & (x8 | (x4 & ~x8)))))) : ((x4 & (x3 ? (x6 & (~x5 | ~x8)) : (~x5 & ~x6))) | (~x4 & ~x5 & ~x6 & x8))))) | (x0 & ~x2 & x3 & x4 & x5 & ~x6 & x8))) | (~x1 & ((~x5 & (x0 ? (x6 ? ((x4 & ((x2 & (x3 ? x7 : (~x7 & x8))) | (x7 & x8 & ~x2 & x3))) | (~x2 & x7 & (x3 ? ~x4 : x8))) : (x4 ? ((~x3 & x7 & ~x8) | (~x7 & (x8 ? x2 : x3))) : (x2 ? (x3 & (~x7 ^ ~x8)) : (~x3 & (~x7 | ~x8))))) : ((x2 & ((x3 & ((x6 & ~x7 & ~x8) | (x4 & x7 & x8))) | (x6 & x7 & ~x8 & ~x3 & x4))) | (~x3 & ((~x6 & ~x7 & x8) | (~x4 & (~x6 | (~x7 & ~x8)))))))) | (x5 & ((x2 & (x3 ? ((x7 & (x0 ? (x4 ? (~x6 & ~x8) : (x6 & x8)) : (x6 & ~x8))) | (~x6 & ~x7 & x8 & ~x0 & ~x4)) : ((x6 & ~x7 & ~x8) | (~x6 & x7 & x0 & ~x4)))) | (x0 & ~x2 & ((~x3 & ~x6 & (x4 ? (~x7 & ~x8) : (x7 & x8))) | (x3 & x4 & x6 & ~x7))))) | (~x2 & (~x0 | (x0 & ~x4 & ~x7 & (x3 ? (x6 & x8) : (~x6 & ~x8))))))) | (x5 & ((x0 & ~x4 & ((~x6 & x7 & x8 & x2 & ~x3) | (x6 & ~x7 & ~x8 & ~x2 & x3))) | (x7 & x8 & x4 & ~x6 & ~x0 & x2 & ~x3)));
  assign z15 = ~x0 & (x1 ? ((x6 & ((~x2 & x5 & (x3 ? (~x4 & ~x7) : (x4 & x7))) | (~x5 & ~x7 & x8 & x2 & ~x3 & ~x4))) | (~x2 & x3 & ((~x4 & x5 & x7) | (~x7 & ~x8 & ~x5 & ~x6)))) : ((~x3 & ((~x4 & (~x6 | (x2 & x6))) | (~x5 & ((~x6 & ~x7 & x8) | (x2 & x4 & (x6 ? (x7 & ~x8) : (x7 | (~x7 & ~x8)))))))) | ~x2 | (x2 & ((x4 & ~x5 & x6 & (~x7 | (x3 & x7))) | (x3 & x5 & ~x6 & (~x8 | (~x7 & x8)))))));
  assign z16 = ~x0 & ((~x7 & ((x6 & ((~x3 & ((~x5 & (x1 ? (x8 & (~x2 ^ ~x4)) : (x2 & x4))) | (~x1 & x2 & ~x4 & x5 & x8))) | (x4 & x5 & ~x8 & x1 & ~x2 & x3))) | (~x1 & ~x6 & ((x2 & ~x8 & (x3 ? ~x4 : (x4 & ~x5))) | (~x3 & ~x5 & x8))))) | (~x2 & (~x1 | (x6 & x7 & ~x8 & x1 & ~x3 & x4))) | (~x1 & ~x3 & ((~x4 & ~x6) | (x2 & (x5 ? (x6 & (x8 ? x7 : ~x4)) : (x4 ? (x7 & (~x6 | (x6 & ~x8))) : x6))))));
  assign z17 = ~x0 & ((~x2 & (~x1 | (x1 & ((x4 & (x3 ? ((x7 & x8 & ~x5 & ~x6) | (~x7 & ~x8 & x5 & x6)) : (x6 & x8 & (~x5 ^ x7)))) | (x6 & ~x7 & ~x8 & ~x3 & ~x4 & x5))))) | (~x1 & ((~x3 & ~x4 & ~x6) | (x2 & ((~x3 & x6 & (x4 ? (x7 & (x5 ^ ~x8)) : (~x5 | (x5 & ~x7)))) | (~x6 & ~x7 & x8 & x3 & ~x4 & x5))))));
  assign z18 = ~x0 & (x1 ? (~x2 & ((x6 & ((~x3 & ~x8 & (x4 ? (~x5 & x7) : (x5 & ~x7))) | (x3 & ~x4 & x5 & ~x7))) | (x3 & ((~x4 & x5 & x7) | (~x5 & ~x6 & ((~x7 & ~x8) | (x4 & x7 & x8))))))) : ((x2 & ((x3 & ((x4 & (x5 ? (~x6 & ~x7) : x6)) | (~x6 & ~x8 & ((x5 & x7) | (~x4 & ~x5 & ~x7))))) | (x6 & x7 & ~x8 & ~x3 & x4 & ~x5))) | ~x2 | (~x3 & ~x4 & ~x5 & (~x6 | (~x7 & ~x8)))));
  assign z00 = 1'b0;
endmodule