module pla__opa ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68;
  assign z00 = ~x00 & ((x01 & (x03 ? (~x04 & ((x02 & (~x05 | x06)) | (~x05 & x06))) : (x05 & (x02 ? ~x04 : (x04 & x06))))) | (x03 & ((x05 & ((~x01 & (x04 | (x02 & x06 & ~x13))) | (x04 & ~x06))) | (~x01 & ~x04 & ~x05 & ~x06))));
  assign z01 = ~x00 & ((~x02 & ((~x01 & (x05 | x06)) | (~x03 & (x04 | x06)))) | (~x01 & (x03 | x04)) | ((~x04 | ~x06) & (x03 | (x01 & x02))) | (x02 & (~x05 | (x03 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 | x09)))) | (x01 & ~x05));
  assign z02 = ~x00 & ((x03 & ((x01 & (x02 ? (x04 & x06 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 | x09)) : (~x04 & ~x06))) | (~x04 & x05 & (~x02 | ~x06 | (~x01 & x13))))) | (~x05 & ((x02 & (~x03 | (~x01 & x06))) | x04 | (x01 & ~x03))) | (~x03 & ((x04 & (~x01 | ~x06)) | (~x02 & ((~x01 & (x05 | x06)) | (~x04 & x06))))) | (~x01 & ~x02 & ~x04 & (x05 | x06)));
  assign z03 = ~x06 & x05 & x04 & x03 & x02 & ~x00 & ~x01;
  assign z04 = ~x06 & x05 & x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z05 = x06 & ~x05 & x04 & x03 & ~x02 & ~x00 & x01;
  assign z06 = ~x06 & ~x05 & x04 & x03 & ~x02 & ~x00 & x01;
  assign z07 = ~x06 & x05 & ~x04 & x03 & x02 & ~x00 & x01;
  assign z08 = x06 & x05 & ~x04 & x03 & x02 & ~x00 & ~x01;
  assign z09 = x06 & x05 & ~x04 & ~x03 & ~x02 & ~x00 & x01;
  assign z10 = ~x06 & ~x05 & ~x04 & ~x03 & x02 & ~x00 & x01;
  assign z11 = ~x16 & ~x15 & ~x14 & ~x12 & ~x09 & x08 & x07 & x06 & x05 & x04 & x03 & x02 & ~x00 & x01;
  assign z12 = ~x16 & ~x15 & ~x14 & ~x12 & ~x09 & x08 & ~x07 & x06 & x05 & x04 & x03 & x02 & ~x00 & x01;
  assign z13 = ~x16 & ~x15 & ~x14 & ~x12 & ~x09 & ~x08 & ~x07 & x06 & x05 & x04 & x03 & x02 & ~x00 & x01;
  assign z14 = ~x00 & x03 & ~x04 & ((x05 & (~x02 | (~x01 & ~x06))) | (~x01 & x06 & (~x02 | ~x05)) | (x01 & ~x02 & ~x06));
  assign z15 = ~x00 & ((~x10 & ((~x03 & ((~x01 & ~x02 & (x05 | x06)) | (x01 & ((x02 & (~x04 | ~x06)) | ~x05 | (~x04 & x06))) | (x04 & ~x06) | (x02 & ~x05))) | (x02 & ((x01 & ~x05) | (x03 & x04 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 | x09)))) | (~x01 & x04))) | (x02 & ((x01 & x05 & (x03 ? ~x06 : ~x04)) | (x03 & x04 & (~x05 | ~x06 | (x07 & ~x08 & x09 & ~x12 & ~x14 & ~x15 & ~x16))))) | (x03 & x04 & (~x01 | (x05 & ~x06) | (~x05 & x06))));
  assign z16 = ~x00 & x10 & ((x01 & ((x02 & ((x03 & x04 & x05 & x06 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 ^ x09)) | (~x04 & ~x05))) | (~x03 & ~x05))) | (~x03 & ((x04 & (~x01 | ~x06)) | (~x02 & ((~x01 & (x05 | x06)) | (~x04 & x06))) | (x02 & ~x05))));
  assign z17 = ~x00 & ((~x03 & ((~x01 & (x04 | (~x02 & x06))) | (~x06 & (x04 | (x01 & x02 & ~x05))) | (~x02 & ~x04 & x06))) | (x01 & ((x04 & ~x05) | (~x04 & ~x06 & ~x02 & x03))) | (~x06 & ((x04 & ~x05) | (x03 & ~x04 & x05))) | (x03 & ~x04 & x05 & (~x01 | ~x02)));
  assign z18 = ~x00 & ((x06 & ((x01 & x05 & (x02 ? (x03 & ~x04) : (~x03 & x04))) | (~x04 & ~x05 & ~x02 & x03))) | (~x04 & ~x05 & ~x01 & x03));
  assign z19 = ~x00 & x03 & ((x01 & ((x02 & ~x04 & ~x05) | (x05 & ~x06 & ~x02 & x04))) | (~x01 & ~x02 & x04 & x05 & x06));
  assign z20 = ~x00 & (x01 ? (~x06 & ((x02 & x03 & x04 & x05) | (~x04 & ~x05 & ~x02 & ~x03))) : (x03 & x04 & x06 & (x02 | ~x05)));
  assign z21 = ~x00 & ((x02 & ((x06 & ((x01 & x03 & x04 & x05 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 | x09)) | (~x03 & ~x04 & ~x05))) | (~x04 & ~x05 & ~x01 & ~x03))) | (~x01 & ~x02 & ~x03 & ~x04 & x05 & ~x06));
  assign z22 = ~x00 & x03 & ((x02 & ((~x01 & x04 & ~x05) | (x05 & ~x06 & x01 & ~x04))) | (x01 & x04 & ~x05 & (x06 | x11)));
  assign z23 = ~x00 & x03 & x04 & ~x05 & ((x02 & (~x01 | ~x06)) | (x01 & ~x02 & x06));
  assign z24 = ~x00 & x01 & x02 & x03 & (x04 ? (~x05 & x06) : (x05 & ~x06));
  assign z25 = ~x00 & ((x05 & ((x03 & ((x01 & x02 & x04 & x06 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 | x09)) | (~x04 & (~x02 | (~x01 & (~x06 | x13)))))) | (~x01 & ~x02 & (~x03 | ~x04)))) | (~x02 & ((x01 & ~x06 & (~x05 | (x03 & ~x04))) | (~x01 & x04 & ~x05) | (x06 & ((~x03 & ~x04) | (~x01 & (~x03 | ~x04)))))) | (~x01 & (x04 ? ~x03 : (~x05 & x06))) | (~x03 & ((x04 & ~x06) | (~x05 & (x01 | x02)))));
  assign z26 = ~x00 & ((x03 & ((~x01 & ((x02 & (x04 | (x05 & x06 & ~x13))) | (x04 & x05) | (~x04 & ~x05 & ~x06))) | (x01 & ((~x05 & x06) | (x02 & (~x04 | ~x05)))) | (x02 & ~x05 & ~x06))) | (x01 & x05 & ((x02 & ~x04) | (x04 & x06 & ~x02 & ~x03))));
  assign z27 = ~x00 & ((x01 & ((~x06 & ((~x02 & (x03 | x04)) | (x04 & x05) | (x02 & ~x03))) | (x02 & ((x03 & x04 & x05 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 | x09)) | (~x04 & (~x03 | (~x05 & x06))))) | (~x03 & (~x05 | (~x04 & x06))))) | (~x01 & ((~x03 & (x04 | (~x02 & x05))) | (~x02 & ((~x04 & x05) | x06 | (x04 & ~x05))) | (x03 & ((~x04 & (x05 | x06)) | (x05 & x06))))) | (x02 & ~x03 & ~x05) | (~x02 & x03 & ~x04 & x05));
  assign z28 = ~x00 & ((x03 & ((x01 & ((x02 & x04 & x05 & ~x08 & ~x12 & ~x14 & ~x15 & ~x16 & (x07 | x09)) | (~x04 & x06) | (~x02 & ~x06))) | (~x02 & (~x04 | (~x01 & ~x05))) | (~x01 & ~x04 & (~x06 | x13)))) | (x01 & ((~x03 & ~x05) | (x05 & ~x06 & x02 & x04))) | (x02 & ~x05 & (~x03 | (~x01 & ~x04))) | (~x01 & ((~x02 & (x06 | (~x03 & x05))) | (x04 & (~x03 | (x05 & x06))))) | (~x03 & ((x04 & ~x06) | (~x02 & (x04 | x06)))));
  assign z29 = ~x00 & x03 & ((x01 & ((x04 & ~x05 & x06) | (x02 & ~x04 & x05 & ~x06))) | (x02 & x04 & ~x05));
  assign z30 = ~x00 & ((x06 & (x01 ? (x02 & ~x04) : (~x02 & ~x03))) | (x02 & ((x01 & ~x04 & (x03 ^ x05)) | (~x01 & (x03 ^ ~x05)) | (x03 & x04 & x05 & ~x08 & x09 & ~x12 & ~x14 & ~x15 & ~x16))) | (~x01 & (x04 | (~x02 & ~x03 & x05))) | (~x02 & ((x04 & ~x05) | (~x03 & (x04 | (x01 & ~x05))))) | (x04 & (~x06 | (~x03 & ~x05))));
  assign z31 = ~x00 & x03 & ((~x02 & ~x04 & ~x05 & (~x01 | ~x06)) | (x01 & x02 & x04 & x05 & x06 & x07 & ~x14 & ~x15 & ~x16 & ~x08 & ~x09 & ~x12));
  assign z32 = ~x00 & ((x04 & ((~x03 & (~x02 | ~x05)) | ~x01 | ~x06 | (x02 & x03 & x05 & ~x12 & ~x14 & ~x15 & ~x16 & ((~x08 & x09) | (x07 & (~x08 | ~x09)))))) | (~x06 & ((x03 & x05 & ~x01 & x02) | (x01 & ~x02 & ~x05))) | (x02 & ((~x01 & ~x03 & ~x05) | (x01 & x03 & ~x04 & x05 & x06))) | (~x03 & ((x01 & ~x05 & (~x02 | x06)) | (~x02 & (x06 | (~x01 & x05))))) | (~x01 & ~x02 & x03 & ~x05));
  assign z33 = ~x00 & x02 & x05 & ((~x03 & ~x04) | (x01 & x03 & x04 & x06 & ~x07 & ~x14 & ~x15 & ~x16 & ~x09 & ~x12));
  assign z34 = ~x00 & ((x06 & ((~x03 & (x02 ? (~x05 & x12) : (x01 ? (x04 & x12) : ~x05))) | (x01 & x02 & x03 & x05 & ((~x04 & x12) | (~x12 & ~x14 & ~x15 & ~x16 & ~x08 & x09 & x04 & ~x07))))) | (~x03 & ((x04 & ~x05) | (~x01 & x12 & ((x02 & ~x05) | (x05 & ~x06 & ~x02 & ~x04))))));
  assign z35 = ~x00 & ((x02 & ((~x01 & ~x03 & ~x05) | (x06 & ((~x03 & ~x05) | (x01 & x03 & x05 & (~x04 | (~x12 & ~x14 & ~x15 & ~x16 & ~x07 & ~x08 & x09))))))) | (~x03 & ((~x01 & (x04 | (~x02 & x05 & ~x06))) | (x04 & (~x02 | ~x05 | ~x06)))));
  assign z36 = ~x00 & x01 & ~x03 & x04 & (~x05 | ~x06);
  assign z37 = ~x00 & x04 & (x01 ? (x06 & ((~x03 & ~x05) | (x09 & ~x12 & ~x14 & ~x15 & ~x16 & x02 & x03 & x05 & ~x07 & ~x08))) : (~x03 & ~x06));
  assign z38 = ~x00 & ((x02 & ((~x01 & ~x03 & ~x05) | (x06 & ((~x03 & ~x05) | (x01 & x03 & x05 & (~x04 | (~x12 & ~x14 & ~x15 & ~x16 & ~x07 & ~x08 & x09))))))) | (~x03 & ((x04 & (~x02 | ~x05 | ~x06)) | (~x01 & (x04 | (~x02 & (x05 | x06)))))));
  assign z39 = ~x00 & ((~x03 & ((~x01 & (x04 | (~x02 & x06))) | (x04 & (~x05 | ~x06)))) | (~x12 & ~x14 & ~x15 & ~x16 & ~x07 & ~x08 & x09 & x04 & x05 & x06 & x01 & x02 & x03));
  assign z40 = ~x00 & x02 & x05 & ((~x03 & ~x04 & ~x06) | (x01 & x03 & x04 & x06 & ~x07 & ~x14 & ~x15 & ~x16 & x08 & ~x09 & ~x12));
  assign z41 = ~x00 & x02 & x05 & ((~x03 & ~x04) | (x01 & x03 & x04 & x06 & ~x07 & ~x14 & ~x15 & ~x16 & x08 & ~x09 & ~x12));
  assign z42 = ~x00 & ((~x03 & ((x02 & ~x04 & ~x05 & (~x01 | x06)) | (x05 & ((~x01 & (~x02 | x04)) | (x04 & (~x02 | ~x06)))))) | (~x04 & x05 & x06 & x01 & x02 & x03));
  assign z43 = x05 & ~x04 & ~x03 & ~x00 & x02;
  assign z44 = ~x00 & ((~x03 & ((~x01 & (x05 | (x02 & ~x04))) | (x02 & ((x05 & ~x06) | (~x04 & (x05 | x06)))) | (~x02 & x04 & x05))) | (x01 & x02 & ~x04 & x05 & x06));
  assign z45 = x05 & ~x04 & ~x03 & x02 & ~x00 & x01;
  assign z46 = ~x00 & x05 & ((x02 & ((x01 & x03 & x04 & x06 & ~x07 & ~x14 & ~x15 & ~x16 & x08 & ~x09 & ~x12) | (~x01 & ~x03 & (~x04 | ~x06)))) | (~x03 & x04 & ~x06));
  assign z47 = ~x00 & x02 & ((x01 & x06 & ((~x03 & ~x04) | (~x14 & ~x15 & ~x16 & ~x09 & ~x12 & x03 & x04 & x05 & ~x07 & x08))) | (~x03 & ((x05 & (~x01 | ~x04)) | (x04 & (~x05 | ~x06)) | (~x01 & (x04 | ~x06)))));
  assign z48 = ~x00 & ((x03 & ((~x01 & (x04 | (x02 & x05 & ~x06))) | (~x02 & ~x05 & (x04 | (x01 & ~x06))) | (x04 & (~x06 | (x02 & x05 & ~x12 & ~x14 & ~x15 & ~x16 & ((x07 & (~x08 | ~x09)) | (~x08 & ~x09))))))) | (x01 & ~x02 & ~x03 & ~x04 & (~x05 | x06)));
  assign z49 = ~x00 & x03 & x04 & (~x01 | ~x06 | (x09 & ~x12 & ~x14 & ~x15 & ~x16 & x02 & x05 & x07 & ~x08));
  assign z50 = ~x00 & x03 & x04 & ((~x05 & (~x01 | ~x06)) | (x01 & x02 & x05 & x06 & x07 & ~x14 & ~x15 & ~x16 & ~x08 & x09 & ~x12));
  assign z51 = ~x00 & x03 & x04 & ((x01 & x02 & x05 & x06 & x07 & ~x14 & ~x15 & ~x16 & ~x08 & x09 & ~x12) | (~x05 & (~x06 | (~x01 & ~x02))));
  assign z52 = ~x00 & x03 & x04 & (~x01 | ~x06 | (x02 & (~x05 | (x07 & ~x08 & x09 & ~x12 & ~x14 & ~x15 & ~x16))));
  assign z53 = ~x05 & ~x04 & x03 & ~x02 & ~x00 & ~x01;
  assign z54 = ~x00 & x03 & ((x01 & x02 & x04 & x05 & x06 & x07 & ~x14 & ~x15 & ~x16 & ~x08 & ~x09 & ~x12) | (~x04 & ((~x02 & (~x01 | ~x05)) | (~x01 & (~x05 | x06)))));
  assign z55 = ~x00 & x03 & (x01 ? ((~x02 & ~x04) | (~x14 & ~x15 & ~x16 & ~x08 & ~x09 & ~x12 & x02 & x04 & x05 & x06 & x07)) : (~x04 & (~x05 | (x02 & x06))));
  assign z56 = ~x00 & x03 & ((x01 & x02 & x04 & x05 & x06 & x07 & ~x14 & ~x15 & ~x16 & ~x08 & ~x09 & ~x12) | (~x04 & ((~x01 & (~x05 | (~x02 & x06))) | (~x02 & (x05 ^ ~x06)))));
  assign z57 = ~x00 & x03 & ~x04 & x12 & (~x02 | (~x01 & ~x05));
  assign z58 = ~x05 & ~x04 & x03 & x02 & ~x00 & x01;
  assign z59 = ~x00 & ~x04 & ((~x01 & ~x03 & ~x06 & (~x02 ^ ~x05)) | (x01 & x02 & x03 & x05 & x06));
  assign z60 = ~x00 & ~x03 & x06 & ((x02 & ~x04 & ~x05) | (x04 & x05 & x01 & ~x02));
  assign z61 = 1'b0;
  assign z62 = 1'b0;
  assign z63 = 1'b0;
  assign z64 = 1'b0;
  assign z65 = 1'b0;
  assign z66 = 1'b0;
  assign z67 = 1'b0;
  assign z68 = 1'b0;
endmodule