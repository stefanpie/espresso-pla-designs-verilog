module pla__signet ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38,
    z0, z1, z2, z3, z4, z5, z6, z7  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38;
  output z0, z1, z2, z3, z4, z5, z6, z7;
  assign z0 = (~x03 & ((~x06 & ((x00 & (x07 ? x01 : x08)) | (x01 & x09) | x22 | (x08 & x11))) | (~x01 & ((x10 & ~x14 & ~x17 & x18) | (x15 & ~x24))) | x27 | (~x14 & x16 & x18))) | (x00 & ((~x01 & ~x02 & x03) | (x04 & x05 & x06))) | ((x18 | x22) & ((~x01 & ~x02 & x03) | (x06 & ~x10))) | (x06 & ((~x01 & ((~x08 & (x26 | (x09 & x10))) | (x04 & x11 & x12 & x13))) | (x11 & (x04 ? (~x12 | ~x13) : ~x25)) | ((x15 | x26) & (~x10 | ~x12)) | (x18 & (x21 | (~x17 & ~x20))) | (x09 & ~x10))) | (x24 & (((x15 | x26) & (x16 | (~x16 & (x17 | (x01 & ~x17))))) | (x01 & (x11 | (~x16 & ~x17 & x18))) | (x18 & (x19 | (~x16 & x17))) | (x19 & ~x23 & x26))) | (x14 & ((x11 & (x23 | (~x01 & ~x08))) | (~x01 & ((~x23 & x26) | (x18 & x19))) | (x18 & (x17 | (x01 & ~x17 & x20))))) | (~x14 & x22 & x23 & ~x24);
  assign z1 = (x00 & ((x02 & x03) | (~x01 & ~x03 & ~x06 & x07))) | (x10 & ((x06 & (((x01 | x08) & (x09 | (x12 & x26))) | (x01 & x12 & x15) | (x22 & x23))) | (((~x03 & x18) | (x24 & x26)) & ((x17 & x33) | (x01 & ~x17 & ~x20 & ~x34))) | ((x16 | (x01 & x33)) & ((x24 & (x15 | x26)) | (~x03 & ~x14 & x18))) | (x15 & x24 & ((x17 & x33) | (x01 & ~x17 & ~x20 & ~x32))) | (~x14 & x16 & x27))) | (x19 & ((x02 & x03 & x22) | (~x01 & x15 & ~x17 & x23 & x24))) | (x03 & ((x02 & (x15 | x18)) | (~x01 & x18 & ~x19) | (x15 & x31))) | (~x01 & ((~x08 & x11 & x24) | (~x03 & x09 & ~x28))) | (x11 & ((x01 & x04 & x06 & x12 & x13) | (~x08 & x24 & x29 & ~x30))) | (x14 & ((x01 & ((~x30 & ((~x08 & (x22 | x27)) | (x18 & x20))) | x15 | (x18 & x20 & x33))) | (x17 & x18 & ~x30))) | (~x06 & x22 & x23) | (~x08 & ~x16 & x24 & x27);
  assign z2 = (x24 & ((~x17 & (x01 ? (~x20 & (x15 | x26)) : (x19 & (x23 ? x26 : x15)))) | ((x15 | x26) & (x16 | (~x33 & (x01 | x17)))) | (x01 & x11))) | (x06 & (((x09 | x26) & (x08 | ~x10)) | (x15 & (~x10 | ~x12)) | (~x10 & (x18 | x22)) | (~x12 & (x26 | (x04 & x11))) | (x04 & ((x00 & x05) | (x11 & ~x13))) | (~x04 & x11 & ~x25))) | (~x03 & ((~x06 & ((x00 & (x07 ? x01 : x08)) | x09 | (x08 & x11))) | (x18 & ((~x14 & (x16 | (x01 & (~x33 | (~x17 & ~x20))))) | (x17 & ~x33))))) | ((x27 | (x22 & ~x23)) & (~x14 | (x14 & (x01 | x08)))) | (x14 & (((x01 | x23) & (x11 | x26)) | (x01 & x18 & ((x20 & ~x33) | (~x17 & ~x20 & x34)))));
  assign z3 = x01 & x18 & ((~x17 & (x14 | (x06 & x10 & ~x16))) | (~x02 & x03 & x31));
  assign z4 = (x18 & ((x01 & ~x17 & x20 & ((~x16 & x24) | (x06 & x10 & x35))) | (x06 & x10 & x17 & x35))) | (x01 & ~x16 & ~x17 & x20 & x24 & (x15 | x26));
  assign z5 = x27 & x24 & x08 & ~x16;
  assign z6 = x27 & x06 & ~x10;
  assign z7 = (x36 & ((x24 & (x15 | x26)) | (~x03 & ~x06 & x18))) | (x37 & x38);
endmodule