module pla__pdc ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39;
  assign z00 = ~x03 & ~x04 & (x00 ? ~x01 : (x01 & ~x02 & ~x05 & (x07 | (~x07 & ((~x11 & ~x12 & ((~x13 & ((~x14 & (x08 ? (~x15 & (~x10 | (~x09 & x10))) : (x15 & (x10 | (x09 & ~x10))))) | (~x08 & x14 & ~x15 & (x10 | (x09 & ~x10))))) | (~x08 & x13 & ~x14 & ~x15 & (x10 | (x09 & ~x10))))) | (~x08 & ~x09 & ~x10))))));
  assign z01 = ~x03 & x04 & (x00 ? ~x01 : (x01 & ~x02 & ~x05 & (x07 | (~x07 & ((~x08 & ~x09 & ~x10) | (~x11 & ~x12 & ((~x08 & x13 & ~x14 & ~x15 & (x10 | (x09 & ~x10))) | (~x13 & ((~x08 & x14 & ~x15 & (x10 | (x09 & ~x10))) | (~x14 & (x08 ? (~x15 & (x09 ^ x10)) : (x15 & (x10 | (x09 & ~x10))))))))))))));
  assign z02 = ~x03 & ~x04 & (x00 ? (~x01 & x05) : (x01 & ~x02 & ~x05 & x06 & (x07 | (~x07 & ((~x11 & ~x12 & ((~x13 & ((~x14 & (x08 ? (~x15 & (~x10 | (~x09 & x10))) : (x15 & (x10 | (x09 & ~x10))))) | (~x08 & x14 & ~x15 & (x10 | (x09 & ~x10))))) | (~x08 & x13 & ~x14 & ~x15 & (x10 | (x09 & ~x10))))) | (~x08 & ~x09 & ~x10))))));
  assign z03 = ~x03 & ((~x00 & ~x02 & ((x06 & (((x09 ^ x10) & ((~x01 & x07 & ((x12 & ((x14 & ((x04 & x05 & x08 & x11 & (x13 ^ x15)) | (~x04 & ~x05 & ~x08 & ~x11 & x13 & ~x15))) | (~x04 & ~x05 & ~x08 & ~x11 & ~x13))) | (~x04 & ~x05 & ~x08 & ~x11 & ~x12 & x14 & ~x15))) | (x01 & x04 & ~x05 & ~x07 & x08 & ~x11 & ~x12 & ~x13 & ~x14 & ~x15))) | (x04 & ((~x11 & ((~x08 & (x01 ? (~x05 & ~x07 & ~x12 & (x10 | (x09 & ~x10)) & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))) : ((x05 & ((~x15 & ((x07 & ((~x10 & ((x09 & x14 & (~x12 | (x12 & x13))) | (~x09 & x12 & ~x13 & ~x14))) | (~x09 & ~x12 & x14))) | (x09 & x10 & x14 & (~x12 | (x12 & x13))))) | (x09 & x12 & ~x13 & ((x10 & (~x14 | (x14 & x15))) | (x07 & ~x10 & ~x14))))) | (x07 & x09 & x12 & ~x13 & x14 & x15 & (~x10 | (~x05 & x10)))))) | (~x01 & ((x05 & ((x08 & ((x07 & (x09 ? ((x12 & ~x13 & ~x14) | (x14 & ~x15 & x10 & ~x12)) : (~x10 & (x12 ? (x13 ? (x14 & ~x15) : ~x14) : (x14 & ~x15))))) | (~x09 & x10 & (x12 ? (x13 ? (x14 & ~x15) : (~x14 | (x14 & x15))) : (x14 & ~x15))))) | (x10 & x12 & ~x13 & x14 & ~x15))) | (~x05 & x07 & x08 & ~x09 & x10 & x12 & ~x13 & x14 & x15))))) | (x01 & ~x05 & (x07 | (~x09 & ~x10 & ~x07 & ~x08))) | (~x01 & x05 & ((x07 & ((x11 & (((x12 ? (~x13 & ~x14) : (x14 & ~x15)) & (~x10 | (x08 & ~x09 & x10))) | (x10 & x12 & ((~x13 & x14 & ~x15) | (x09 & ((~x13 & ~x14) | (~x08 & x14 & (x13 ^ x15)))))))) | (x12 & ((x14 & (((x13 ^ x15) & (x08 ? (x09 & x10) : ~x09)) | (~x10 & ~x13 & ~x15))) | (~x08 & ~x09 & x10 & ~x13 & ~x14))))) | (~x10 & x11 & x12 & x14 & (x13 ^ x15) & (~x08 ^ ~x09)))))) | (~x01 & ~x04 & ~x05 & (x07 ? (~x09 & ~x10 & (x08 ^ x11) & (x12 ? (~x13 | (x13 & x14 & ~x15)) : (x14 & ~x15))) : ((x14 & ~x15) | (x12 & ~x13 & (~x14 | (x14 & x15)))))))) | (~x01 & ((~x06 & (x04 ? ((~x15 & (x07 ? ((~x10 & (x12 ? ((~x08 & (x05 ? ((~x11 & x13 & x14) | (~x09 & ~x13 & ~x14)) : ((~x11 & (x09 ? (x14 | (~x13 & ~x14)) : (x13 & x14))) | (~x09 & x11 & ~x13)))) | (~x11 & ((~x05 & ((x08 & x09 & (~x13 | (x13 & x14))) | (~x09 & ~x13))) | (x08 & ~x09 & x13 & x14))) | (x11 & x14 & (x13 | (~x05 & x09 & ~x13)))) : (x14 & (x11 ? (x09 | (~x08 & ~x09)) : ((x08 & (x09 ? ~x05 : ~x13)) | (~x08 & (~x13 | (x09 & x13))) | (~x09 & x13)))))) | (x14 & ((x12 & (x05 ? (~x13 | (x10 & x13)) : ((x08 & x11 & (x13 ? x10 : ~x09)) | (x10 & ~x11)))) | (x10 & ((~x11 & ~x12) | (~x05 & x11 & (~x08 | (x08 & x09 & ~x12))))) | (x08 & ~x09 & x11 & ~x12))) | (~x05 & x08 & x09 & x10 & x11 & x12 & ~x13)) : (x14 & (~x05 | (x05 & ~x11 & ~x12 & ~x13 & (~x08 ^ ~x09)))))) | (x12 & ~x13 & ((~x05 & (x07 ? ((~x14 & (x11 ? ((x08 & (~x09 | (x09 & x10 & x15))) | (x09 & ~x10) | (~x08 & x10)) : (x10 | (~x09 & ~x10 & x15)))) | (~x10 & ~x11 & x15 & (x09 | (~x08 & ~x09 & x14)))) : (~x14 | (x14 & x15)))) | (x07 & (x10 ? (x14 ? x15 : x05) : ((x15 & ((~x08 & ((x05 & ~x11 & x14) | (~x09 & x11 & ~x14))) | (x11 & x14))) | (x05 & ~x14 & (x09 | (x08 & ~x09))))))))) : (x05 & ((~x11 & (x07 ? (~x08 ^ ~x09) : ((~x10 & ((x14 & ~x15 & (~x12 | (x12 & x13)) & (~x08 | (x08 & x09))) | (x12 & ~x13 & (~x08 | (x08 & ~x09))))) | (x08 & (x09 ? (x12 & ~x13) : (x14 & ~x15 & (~x12 | (x12 & x13)))))))) | (~x07 & ((x14 & ~x15 & (~x12 | (x12 & x13)) & (x10 ? (x09 | (~x09 & (~x08 | (x08 & x11)))) : x11)) | (x12 & ~x13 & (x10 ? (~x08 | (x08 & (~x09 | (x09 & x11)))) : x11)))))))) | (x04 & x07 & ((x05 & (x08 ? (x09 & x14 & ((~x10 & ~x11 & (x12 ? (x13 ^ x15) : ~x15)) | (x10 & x11 & ~x12 & ~x15))) : ((~x09 & ~x10 & ~x11 & ~x14 & x15 & x12 & ~x13) | (~x12 & x14 & ~x15 & x10 & x11)))) | (x08 & ~x09 & ~x10 & ~x11 & x14 & x15 & x12 & ~x13))))))) | (x00 & ~x01 & x04 & x05));
  assign z04 = ~x00 & ~x01 & ~x02 & ~x03 & (x04 ? (((~x08 ^ ~x09) & ((x06 & ((x05 & (x11 ? (((~x10 | (x07 & x10)) & (x12 ? (x13 & (~x14 | (x14 & ~x15))) : (x14 & x15))) | (~x13 & x14 & x15 & ~x10 & x12)) : (x14 & ((x12 & (x13 ^ x15) & (x10 | (x07 & ~x10))) | (x07 & ~x10 & ~x12 & x15))))) | (x07 & x11 & x12 & ~x13 & x14 & x15 & (x10 | (~x05 & ~x10))))) | (x05 & ~x06 & ~x07 & x11 & x14 & ~x15 & ~x12 & ~x13))) | (x12 & ((~x06 & ((~x05 & (x07 ? ((~x11 & (x10 ? (x13 & ((x14 & (~x15 | (x09 & x15))) | (~x08 & ~x09 & x15))) : ((x15 & (x08 ? (x09 ? (x13 | (~x13 & x14)) : (x13 & ~x14)) : (x13 | (~x09 & ~x13 & x14)))) | (x13 & (x08 ? (~x09 & x14) : (~x15 & (~x14 | (~x09 & x14)))))))) | (x13 & ((x10 & (x08 ? ((x11 & ((x14 & ~x15) | (x09 & (x15 | (~x14 & ~x15))))) | (~x09 & x14 & x15)) : (x11 & x14))) | (x14 & x15 & ~x10 & x11)))) : (x13 | (~x13 & x14 & x15)))) | (x07 & (x13 ? ((~x11 & ((~x14 & ((x05 & x15 & (x08 ? ~x10 : ~x09)) | (x09 & x10) | (~x09 & ~x15 & (x08 ^ x10)))) | (~x10 & ~x15 & ((x09 & (x08 | (~x08 & x14))) | (x05 & ~x09 & x14))))) | (x14 & ((x05 & (x15 | (x10 & ~x15))) | (~x10 & x11 & ~x15))) | (~x14 & (x10 ? (x08 ? ~x09 : x11) : x11))) : (x14 & x15 & (x10 | (~x10 & (x11 | (~x11 & (x09 ? ~x08 : x05)))))))))) | (x05 & ((x07 & ((x06 & (x13 ? ((x08 & ((x09 & (x14 ? ~x15 : ~x10)) | (~x09 & ~x10 & ~x11 & ~x14))) | (x10 & (x11 ? (x14 & x15) : ~x14)) | (~x11 & x15 & (x14 | (~x10 & ~x14 & ~x08 & ~x09))) | (~x08 & ~x09 & (x14 ? ~x15 : x11))) : (x14 & x15 & (x08 ? (x09 & (x10 | (~x10 & x11))) : ~x09)))) | (x09 & ((x08 & ((x10 & x11 & x13 & ~x14) | (~x13 & x14 & x15 & ~x10 & ~x11))) | (~x08 & ~x10 & ~x11 & x13 & ~x14))) | (~x08 & ~x09 & ~x10 & ~x14 & ~x15 & ~x11 & x13))) | (x06 & ~x10 & x11 & x13 & x14 & x15))))) | (x14 & x15 & ((x07 & ((~x12 & ((~x11 & ((~x06 & ((~x10 & ((~x08 & (~x13 | (x09 & x13))) | (~x05 & (x09 ? x08 : x13)))) | (x09 & x10) | (~x09 & (x08 ? x05 : x10)))) | (x05 & ((x06 & (x10 | (~x08 & ~x09 & ~x10 & ~x13))) | (~x10 & (x08 ? x09 : (~x09 & x13))))))) | (x11 & (x05 ? (~x06 | (x06 & (x08 ^ ~x09))) : (~x06 & (~x10 | (x10 & (~x08 | (x08 & x09))))))) | (x08 & ~x09 & x10 & ~x05 & ~x06))) | (~x05 & ~x06 & x08 & ~x09 & ~x10 & ~x11 & ~x13))) | (~x05 & ~x06 & ~x07 & ~x12)))) : (x05 ? (~x06 & ((x11 & (x07 ? (~x08 ^ ~x09) : ((x14 & x15 & (~x10 | (x08 & ~x09 & x10)) & (~x12 | (x12 & ~x13))) | (x12 & x13 & (~x10 | (x08 & x09 & x10)))))) | (~x07 & ((x14 & x15 & (~x12 | (x12 & ~x13)) & ((~x11 & (x08 ? (~x09 | (x09 & ~x10)) : ~x10)) | (x10 & (x09 | (~x08 & ~x09))))) | (x12 & x13 & (((~x08 | (x08 & ~x09)) & (x10 | (~x10 & ~x11))) | (x08 & x09 & ~x11))))))) : (x06 & (x12 ? (x13 | (~x13 & x14 & x15)) : (x14 & x15)) & (~x07 | (x07 & ((x08 & ~x09 & ~x10 & ~x11) | (~x08 & (x09 ? (~x10 & ~x11) : (~x10 ^ ~x11)))))))));
  assign z05 = ~x00 & ~x01 & ~x02 & ~x03 & ((((~x12 & (x15 ? ~x14 : x13)) | (~x13 & (x14 ? ~x15 : x12))) & ((~x06 & (x04 ? (~x05 & (~x07 | (x07 & x11 & (x10 ? ~x08 : x09)))) : (x05 & ~x07 & (x08 ? (~x09 & x10) : (x10 | (~x10 & x11)))))) | (~x04 & ~x05 & x06 & ~x07))) | ((~x08 ^ ~x09) & ((~x11 & (x05 ? ((~x06 & ((~x04 & x07) | (~x13 & x14 & ~x15 & x04 & ~x07 & ~x12))) | (x04 & x06 & ((x14 & (x12 ? ((x13 ^ x15) & (x10 | (x07 & ~x10))) : ((x07 & ~x10 & x13 & x15) | (~x07 & x10 & ~x15)))) | (x12 & ~x14 & ((x07 & ~x10 & (~x13 | (x13 & x15))) | (x10 & ~x13)))))) : (x06 & x07 & ((~x10 & ((x14 & x15 & x12 & ~x13) | (~x04 & ((~x13 & (x15 ? ~x14 : x12)) | (~x12 & x14 & ~x15) | (x13 & (x12 ? (~x14 ^ ~x15) : (~x14 | (x14 & x15)))))))) | (~x13 & x14 & x15 & x04 & x10 & x12))))) | (x04 & x05 & x06 & x11 & ((x12 & ((x14 & (x13 ^ x15) & (~x10 | (x07 & x10))) | (~x14 & x15 & ~x10 & x13))) | (x13 & x14 & x15 & ~x10 & ~x12))))) | ((~x14 ^ ~x15) & ((x12 & x13 & (x04 ? ((x07 & ~x10 & ~x11 & (x05 ? (x08 ? x09 : ~x06) : (~x06 & (x08 ^ ~x09)))) | (~x05 & ~x06 & ~x07)) : ((~x09 & ((~x08 & ((~x05 & x06 & x07 & (~x10 ^ ~x11)) | (x05 & ~x06 & ~x07 & x10))) | (x05 & ~x06 & ~x07 & x08 & (~x11 | (x10 & x11))))) | (~x07 & (x05 ? (~x06 & ((x09 & (x10 | (x08 & ~x10 & ~x11))) | (~x10 & (x11 | (~x08 & ~x11))))) : x06))))) | (x04 & x07 & ~x10 & ~x11 & ~x12 & ~x13 & (x05 ? (~x08 | (x08 & (x09 | (x06 & ~x09)))) : (~x06 & ~x08))))) | ((~x12 ^ ~x13) & ((x14 & x15 & (x04 ? ((x07 & ~x10 & ~x11 & (x05 ? (x08 ? x09 : ~x06) : (~x06 & (x08 ^ ~x09)))) | (~x05 & ~x06 & ~x07)) : ((~x09 & ((~x08 & ((~x05 & x06 & x07 & (~x10 ^ ~x11)) | (x05 & ~x06 & ~x07 & x10))) | (x05 & ~x06 & ~x07 & x08 & (~x11 | (x10 & x11))))) | (~x07 & (x05 ? (~x06 & ((x09 & (x10 | (x08 & ~x10 & ~x11))) | (~x10 & (x11 | (~x08 & ~x11))))) : x06))))) | (x04 & ~x05 & ~x06 & x07 & ~x08 & x09 & ~x10 & ~x11 & ~x14 & ~x15))) | (~x06 & (x04 ? (x07 & (((~x14 | (x14 & ~x15)) & ((~x05 & ~x08 & ~x09 & ~x11 & ~x12 & x13) | (x05 & x12 & ~x13))) | (((x11 & ~x14 & x15) | (x10 & x14 & ~x15)) & ((x12 & x13) | (x05 & ~x12 & ~x13))) | (~x11 & ((x15 & (x09 ? ((~x05 & ((~x10 & (x08 ? (~x13 & ~x14) : (x13 ? ~x14 : x12))) | (x10 & ~x12 & x13 & ~x14))) | (x10 & (x12 ? (x13 & ~x14) : (x13 ^ ~x14)))) : (x12 ? ((x08 & ((x13 & ~x14) | (~x10 & ~x13 & x14))) | (~x14 & ((~x08 & x10 & x13) | (~x05 & ~x10 & ~x13)))) : ((x13 ^ ~x14) & (x08 | (~x08 & x10)))))) | (~x05 & ((x09 & ((~x10 & ((x14 & (x08 ? (~x12 & ~x15) : (x12 ? ~x15 : x13))) | (x08 & (x12 ? (~x13 & ~x15) : (x13 & ~x14))))) | (x13 & ~x15 & x10 & ~x12))) | (~x13 & ((x10 & (x14 ? ~x15 : x12)) | (~x09 & ~x10 & x12 & ~x15))))) | (x08 & ~x09 & ~x10 & x14 & ~x15 & (~x12 ^ x13)))) | (x11 & ((~x05 & (((x08 ? (x09 & x10) : (~x09 & ~x10)) & ((~x13 & (x15 ? ~x14 : x12)) | (~x12 & (x14 ? ~x15 : x13)))) | (x08 & ~x09 & ~x13 & (x14 ? ~x15 : (x12 | (~x12 & x15)))))) | (x14 & ((~x10 & x12 & (x13 ^ x15)) | (~x12 & x13 & x15))))) | (x10 & x12 & ~x13 & x14 & x15) | (~x05 & x08 & ~x09 & ~x12 & x13 & (~x15 | (~x14 & x15))))) : (x05 & ~x07 & ((~x10 & (((x08 ? (x11 | (~x09 & ~x11)) : ~x11) & ((~x12 & x14 & ~x15) | (~x13 & (x15 ? ~x14 : x12)))) | (~x12 & x13 & ~x14 & (x11 ? x08 : (~x09 | (~x08 & x09)))))) | (x08 & x09 & (~x11 | (x10 & x11)) & ((~x13 & (x15 ? ~x14 : x12)) | (~x12 & (x14 ? ~x15 : x13)))))))) | (x07 & ((x06 & (x04 ? (x05 & (x14 ? ((x10 & ((x08 & ((x09 & x12 & (x13 ^ x15)) | (~x12 & x13 & x15 & ~x09 & x11))) | (x11 & ((~x13 & ~x15) | (x13 & x15 & ~x08 & ~x12))) | (~x11 & ~x12 & (x13 ^ ~x15)))) | (x13 & (x08 ? (x09 & x11 & ((~x12 & x15) | (~x10 & x12 & ~x15))) : (~x09 & ((x12 & ~x15) | (~x10 & ~x12 & x15))))) | (x12 & ~x13 & ((~x08 & ~x09 & x15) | (~x10 & (~x15 | (x08 & x09 & x11 & x15)))))) : (x12 ? ((x08 & ((x09 & (x11 ? (x13 & x15) : ~x13)) | (~x09 & x10 & x11 & x13 & x15))) | (~x08 & ((~x09 & ((~x11 & ~x13) | (~x10 & x13 & x15))) | (x10 & x11 & x13 & x15))) | (x11 & ~x13) | (x10 & ~x11 & x13 & x15)) : (~x13 & x15 & (x10 | (~x10 & x11)))))) : (~x05 & ~x08 & ~x09 & (~x10 ^ ~x11) & ((~x13 & (x15 ? ~x14 : x12)) | (~x12 & (x14 ? ~x15 : x13)))))) | (x04 & x05 & ~x12 & ((x13 & (~x15 | (~x14 & x15))) | (~x13 & x14 & ~x15 & ~x10 & x11))))) | (x04 & x05 & x06 & x10 & ~x13 & x14 & ~x15 & ~x11 & x12));
  assign z06 = x03 & ~x00 & ~x01;
  assign z07 = ~x03 & ~x04 & ~x05 & (x00 ? ~x01 : (x01 & ~x02 & ~x06 & (x07 | (~x07 & ((~x11 & ~x12 & ((~x13 & ((~x14 & (x08 ? (~x15 & (~x10 | (~x09 & x10))) : (x15 & (x10 | (x09 & ~x10))))) | (~x08 & x14 & ~x15 & (x10 | (x09 & ~x10))))) | (~x08 & x13 & ~x14 & ~x15 & (x10 | (x09 & ~x10))))) | (~x08 & ~x09 & ~x10))))));
  assign z08 = ~x03 & ((~x00 & ~x02 & ((~x11 & ((~x05 & ((x04 & ~x06 & ((~x14 & ((~x08 & ((~x12 & ((x13 & ((~x15 & ((x01 & ~x07 & (x10 | (x09 & ~x10))) | (x09 & ~x10 & ~x01 & x07))) | (~x01 & x07 & ~x09))) | (x01 & ~x07 & ~x13 & x15 & (x10 | (x09 & ~x10))))) | (~x01 & x07 & x15 & (x09 ? (~x10 & x13) : (x12 & (~x13 | (~x10 & x13))))))) | (x08 & ((~x12 & ((x01 & ~x07 & ~x13 & ~x15 & (x09 ^ x10)) | (~x01 & x07 & x09 & ~x10 & x13))) | (~x01 & x07 & x09 & ~x10 & x12 & x13 & x15))) | (~x01 & x07 & x09 & x10 & ~x12 & x13 & x15))) | (~x12 & ((x14 & ((~x01 & x07 & x09 & ~x10 & x13) | (~x08 & ((~x15 & ((x01 & ~x07 & ~x13 & (x10 | (x09 & ~x10))) | (~x09 & x13 & ~x01 & x07))) | (~x10 & x13 & x15 & ~x01 & x07 & ~x09))))) | (~x01 & x07 & x09 & x10 & x13 & ~x15))))) | (~x01 & ~x04 & x06 & x07 & (x13 ? (~x12 | (x12 & ~x14 & x15)) : (~x14 & x15)) & (x08 ? (~x09 & ~x10) : (x09 ^ x10))))) | (~x01 & ((x05 & (x04 ? ((x07 & (x13 ? ((x15 & (x12 ^ x14) & (x10 ? x06 : ((x08 & x09) | (~x06 & ~x08) | (x06 & (~x08 ^ ~x09))))) | (~x12 & ~x15 & ((x14 & ((~x08 & ~x09 & ~x10) | (x06 & x08 & x09))) | (x06 & (x10 ? ~x14 : (x08 ? (~x09 | (x09 & ~x14)) : (x09 | (~x09 & ~x14)))))))) : (~x14 & x15 & ((x12 & ((~x08 & ~x09) | (x06 & x08 & x09))) | (x06 & (x10 ? ~x12 : (x08 ? (~x09 | (x09 & ~x12)) : (x09 | (~x09 & ~x12))))))))) | (x06 & x10 & (~x08 ^ ~x09) & ((~x14 & x15 & x12 & ~x13) | (x14 & ~x15 & ~x12 & x13)))) : (~x06 & ~x07 & ((~x10 & ((~x14 & x15 & (~x08 | (x08 & x09)) & (~x13 | (x12 & x13))) | (~x12 & x13 & (~x09 | (~x08 & x09))))) | (x08 & (x09 ? (~x12 & x13) : (~x14 & x15 & (~x13 | (x12 & x13))))))))) | (x04 & ~x06 & x07 & x15 & (x13 ? ((x12 ^ x14) & (x09 ? x10 : (x08 | (~x08 & x10)))) : (~x14 & (x10 ? (x09 | (~x08 & ~x09 & ~x12)) : (x08 ? x09 : (~x12 | (x09 & x12))))))))))) | (x04 & ((~x06 & ((~x05 & (x01 ? (x07 | (~x09 & ~x10 & ~x07 & ~x08)) : (x07 ? ((x08 & ~x09 & ~x12 & x13 & (~x15 | (~x14 & x15))) | (x11 & ((x13 & (x12 ? (~x14 & x15 & (~x10 | (x08 & x10))) : ((x09 & ((x08 & x10 & (~x14 | (x14 & ~x15))) | (~x10 & (~x15 | (~x14 & x15))))) | (~x08 & ((x10 & ~x15) | (~x09 & ~x10 & ~x14)))))) | (x10 & ~x14 & x15 & (~x08 | (x08 & x09 & ~x13)))))) : ((~x14 & x15) | (~x12 & x13 & (~x15 | (x14 & x15))))))) | (~x01 & x07 & ((~x09 & ((~x10 & ((~x12 & x13 & ~x15 & ((~x08 & x11 & x14) | (x05 & (x08 | (~x08 & ~x14))))) | (~x08 & x11 & ~x13 & ~x14 & x15))) | (~x14 & x15 & x08 & ~x13))) | (x09 & ~x10 & ((~x14 & x15 & x11 & ~x13) | (x13 & ~x15 & x05 & ~x12))) | (x13 & ((x05 & ((~x14 & x15 & x11 & x12) | (x10 & ~x12 & ~x15))) | (x14 & x15 & x11 & ~x12))))))) | (~x01 & x05 & ((x06 & ((x11 & ((x07 & (((~x10 | (x08 & ~x09 & x10)) & ((~x13 & ~x14 & x15) | (~x12 & x13 & ~x15))) | (x13 & ((x10 & ((x15 & (~x08 | (x08 & ~x09)) & (x12 ^ x14)) | (~x12 & ~x15 & (x09 | (~x08 & ~x09 & ~x14))))) | (x08 & x09 & x15 & (x12 ^ x14)))))) | (~x10 & x13 & x15 & (~x08 ^ ~x09) & (x12 ^ x14)))) | (x07 & ~x08 & ~x09 & x13 & ((x14 & ~x15 & x10 & ~x12) | (~x10 & x15 & (x12 ^ x14)))))) | (x07 & ~x14 & x15 & ((~x12 & x13) | (x10 & x11 & ~x13 & (~x08 | (x08 & x09))))))))) | (~x01 & ~x04 & ((x11 & ((~x10 & (x13 ? (~x12 | (x12 & ~x14 & x15)) : (~x14 & x15)) & ((x05 & ~x06 & ~x07) | (~x05 & x06 & x07 & ~x08 & ~x09))) | (x05 & ~x06 & ~x07 & x08 & x10 & (x09 ? (~x12 & x13) : (~x14 & x15 & (~x13 | (x12 & x13))))))) | (~x07 & (x05 ? (~x06 & x10 & ((~x14 & x15 & (x09 | (~x08 & ~x09)) & (~x13 | (x12 & x13))) | (~x12 & x13 & (~x08 | (x08 & ~x09))))) : (x06 & ((~x14 & x15) | (~x12 & x13 & (~x15 | (x14 & x15))))))))))) | (x00 & ~x01 & x04 & ~x05));
  assign z09 = ~x00 & ~x01 & ~x02 & ~x03 & ((x07 & ((~x13 & ((~x12 & (((x15 | (x14 & ~x15)) & ((x06 & ((~x10 & ((~x11 & (~x08 ^ ~x09) & (x04 ^ ~x05)) | (~x04 & ~x05 & ~x08 & ~x09 & x11))) | (~x09 & x10 & ((x08 & x11 & x04 & x05) | (~x04 & ~x05 & ~x08 & ~x11))))) | (x04 & ~x06 & x11 & ((x09 & ~x10) | (~x05 & x10 & (~x08 | (x08 & x09))))))) | (x04 & ((x05 & ((x08 & ((~x06 & ~x09 & (x15 | (~x10 & x14 & ~x15))) | (x09 & (x10 ? ((x11 & x15) | (x06 & x14 & ~x15)) : ((x06 & x15 & (x14 | (~x11 & ~x14))) | (~x11 & x14 & ~x15)))))) | (~x08 & ((x14 & ((~x09 & ~x10 & x15) | (x06 & ~x15 & (x11 ? x10 : ~x09)))) | (x15 & ((x10 & x11) | (~x09 & ~x10 & ~x11 & ~x14))))) | (x10 & (x06 ? (~x11 & x15) : (x14 & ~x15))) | (~x14 & ~x15) | (x06 & ~x10 & x11 & (~x14 ^ ~x15)))) | (~x06 & ((~x05 & ((~x10 & ((~x08 & ((~x09 & x14 & x15) | (~x11 & ~x14 & ~x15))) | (x09 & ~x15 & ((x11 & ~x14) | (x08 & ~x11 & x14))) | (~x09 & ((x08 & (x11 ? x15 : x14)) | (~x11 & ~x14 & x15))))) | (x10 & ((x08 & ~x09 & (x15 | (~x14 & ~x15))) | (~x11 & ~x15 & (x14 | (x09 & ~x14))))) | (x08 & ~x09 & x11 & x14 & ~x15))) | (~x08 & ((~x09 & (x10 ? (~x11 & x15) : (x11 & (~x14 ^ ~x15)))) | (x14 & ~x15 & ~x10 & ~x11))) | (x09 & ~x11 & x15))))))) | (x04 & ~x14 & ~x15 & ((x12 & ((~x06 & ((x05 & (x10 | (x08 & ~x09 & ~x10))) | (~x05 & x10 & (~x11 | (x08 & x11))) | (~x10 & ((x09 & x11) | (~x08 & (~x11 | (~x09 & x11))))))) | (x05 & x06 & (x11 | (~x11 & (x08 ? (x09 | (~x09 & ~x10)) : (~x09 | (x09 & ~x10)))))))) | (~x05 & ~x06 & ((x08 & ~x09 & ~x10 & ~x11) | (~x08 & x10 & x11))))))) | (~x14 & ~x15 & ((~x09 & ((~x08 & ((x06 & (x04 ? (x05 & x13 & ((x11 & (x12 | (x10 & ~x12))) | (~x10 & ~x11 & ~x12))) : (~x05 & (~x10 ^ ~x11)))) | (x04 & ((~x11 & ((x13 & ((x05 & (x12 ? ~x10 : ~x06)) | (~x06 & x10 & x12))) | (x10 & ~x12 & ~x05 & ~x06))) | (~x05 & ~x06 & ~x10 & x12 & x13))))) | (x04 & ((x08 & ((x13 & ((x05 & x06 & (~x10 ^ x11)) | (~x06 & (x10 | (~x10 & ~x11 & x12))))) | (~x05 & ~x06 & ~x10 & x11 & x12))) | (~x05 & ~x06 & ~x10 & ~x12 & (x11 | (~x11 & x13))))) | (x08 & ~x10 & ~x11 & ~x04 & ~x05 & x06))) | (x04 & ((x09 & ((x13 & ((x08 & ((x05 & ((x10 & x11) | (x06 & ~x10 & (x12 | (~x11 & ~x12))))) | (~x05 & ~x06 & x10 & x11 & x12))) | (~x08 & ((x05 & ((~x10 & ~x11) | (x06 & x10 & x11))) | (~x10 & ~x11 & ~x05 & ~x06))) | (~x06 & ((x10 & ~x11) | (~x05 & ~x10 & x11))))) | (~x06 & x08 & ((~x10 & ~x11 & x12) | (~x05 & ~x12 & (~x10 ^ x11)))))) | (x13 & ((x05 & (x06 ? (x10 ? ~x11 : (x11 & ~x12)) : (~x10 & (x11 | (x08 & ~x11 & ~x12))))) | (x10 & x11 & ~x06 & ~x08))))) | (~x04 & ~x05 & x06 & ~x08 & x09 & ~x10 & ~x11))))) | (x05 & (x04 ? (x06 & (~x08 ^ ~x09) & ((~x13 & ((x10 & ~x11 & ~x15 & (x12 ^ x14)) | (~x10 & x11 & ~x12 & x14 & x15))) | (x13 & ~x14 & ~x15 & ~x10 & x11 & x12))) : (~x06 & ~x07 & ((~x12 & ~x13 & (x15 | (x14 & ~x15)) & ((~x08 & (x10 ? ~x09 : ~x11)) | (x09 & (x10 | (x08 & ~x10 & ~x11))) | (~x10 & x11) | (x08 & ~x09 & (~x11 | (x10 & x11))))) | (~x14 & ~x15 & (((~x08 | (x08 & ~x09)) & (x10 | (~x10 & ~x11))) | (~x10 & x11) | (x08 & x09 & (~x11 | (x10 & x11))))))))) | (~x05 & ~x07 & (x04 ^ x06) & ((~x14 & ~x15) | (~x12 & ~x13 & (x15 | (x14 & ~x15))))));
  assign z10 = ~x00 & ~x01 & ~x02 & ~x03 & x04 & x05 & ((~x13 & ((~x12 & (x06 ? (x07 & (x15 | (~x14 & ~x15))) : (~x07 & x14 & ~x15 & (~x08 ^ ~x09)))) | (x06 & x07 & x12 & (~x14 | (x14 & x15))))) | (x06 & x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))))));
  assign z11 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x06 & x07 & ((x08 & ~x09 & ~x10 & ~x11) | (~x08 & (x09 ? (~x10 & ~x11) : (~x10 ^ ~x11))));
  assign z12 = ~x00 & ~x01 & ~x02 & ~x03 & x04 & ~x05 & ~x06 & ~x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))));
  assign z13 = ~x00 & ~x01 & ~x02 & ~x03 & x04 & ~x05 & ~x06 & x07 & ((~x10 & ((~x15 & ((x08 & ((~x09 & x11 & ~x14) | (x09 & ~x11 & ~x12 & ~x13 & x14))) | (x09 & ((x11 & (~x14 | (x12 & ~x13 & x14))) | (~x08 & ~x11 & ((x13 & ~x14) | (x12 & (x14 | (~x13 & ~x14))))))) | (~x08 & ((~x11 & ((~x12 & ~x13) | (~x09 & x12 & x13 & x14))) | (~x09 & x12 & (~x13 | (x13 & ~x14))))))) | (x15 & ((x11 & ((~x14 & ((x08 & (~x13 | (x12 & x13))) | (x09 & ~x12 & x13) | (~x08 & x12))) | (x12 & ~x13 & x14) | (~x08 & ~x12 & (x13 ? x14 : x09)))) | (~x11 & ((x09 & (~x08 | (x13 & x14 & x08 & ~x12))) | (~x08 & ~x09 & ((~x13 & (~x14 | (x12 & x14))) | (~x12 & x13 & x14))))) | (~x08 & ~x09 & ~x12 & ~x13 & x14))) | (~x09 & ((~x11 & ((x08 & (~x13 | (x12 & x13 & x14))) | (x13 & ~x14 & ~x08 & ~x12))) | (~x08 & x11 & ~x12 & ~x14))) | (x08 & ((x09 & ~x11 & (x12 | (~x12 & ~x14))) | (x11 & ~x12 & x14))) | (x13 & x14 & x11 & x12))) | (x10 & ((x08 & ((~x14 & (x09 ? (x11 ? (~x12 | (x12 & (x13 ^ x15))) : (x15 ? ~x13 : x12)) : ((x11 & x13 & (~x15 | (x12 & x15))) | (~x13 & (x12 | (~x12 & ~x15)))))) | (x15 & ((x11 & ((~x12 & x13 & x14) | (x09 & (x12 ? x13 : (~x13 & x14))))) | (~x09 & (x12 ? (x13 & x14) : ~x13)))) | (~x15 & ((x12 & x13 & x14) | (x11 & ((~x12 & x14) | (x09 & x12 & ~x13))))))) | (~x11 & ((x09 & ((x13 & x15) | (~x12 & ~x14 & ~x15))) | (~x13 & x14 & ~x15) | (~x08 & ((~x09 & ~x12 & (~x14 | (x14 & x15))) | (x12 & x13 & ~x15))))) | (x14 & x15 & x12 & ~x13) | (~x08 & ((x12 & ((~x13 & ~x14) | (x11 & x14 & ~x15))) | (x11 & ((x13 & (x15 | (~x14 & ~x15))) | (~x12 & ~x13 & (x15 ? ~x09 : ~x14)))) | (~x13 & x15 & x09 & ~x12))))) | (x08 & ((~x11 & ((~x12 & ((x14 & (x09 ? (x13 ^ x15) : (x13 & x15))) | (~x09 & x13 & ~x15))) | (~x09 & x12 & x13 & ~x14))) | (~x09 & ((~x14 & x15 & ~x12 & x13) | (~x13 & x14 & ~x15 & x11 & x12))))) | (~x08 & ((~x11 & x13 & ((~x12 & x14 & ~x15) | (~x09 & x12 & x15))) | (x14 & ~x15 & x11 & ~x12))));
  assign z14 = x00 & ~x01;
  assign z15 = x00 ? (~x01 & ~x02) : x02;
  assign z16 = ~x00 & ~x01 & ~x02 & ~x03 & x08 & ((x05 & (((~x11 | (x10 & x11)) & ((~x04 & ~x06 & ~x07 & x09) | (x04 & x06 & x07 & x12 & x13 & x15))) | (x04 & ((x06 & ((~x09 & (x10 ? ((x14 & ((~x15 & (~x12 | (x12 & x13)) & (~x11 | (x07 & x11))) | (~x13 & x15 & ~x11 & x12))) | (~x13 & ~x14 & ~x11 & x12)) : ((x11 & ((~x07 & (x12 ? (x13 & ~x14) : (x14 & x15))) | (x12 & x14 & (x13 ^ x15)))) | (x07 & ~x11 & ((x12 & (x13 ? (x14 & ~x15) : ~x14)) | (~x15 & (x14 ? ~x12 : x13))))))) | (x07 & ((x14 & ((~x15 & ((x10 & ((x09 & ~x12) | (x11 & x12 & ~x13))) | (x09 & ((x12 & x13) | (~x10 & ~x11 & ~x12 & ~x13))) | (~x10 & x12 & ~x13))) | (~x13 & x15 & x09 & x12))) | (~x12 & x13 & x15) | (x12 & ~x14 & ((x11 & (~x13 | (~x10 & x13 & x15))) | (x09 & ~x11 & ~x13))))) | (x12 & x14 & ((~x10 & x11 & x13 & x15) | (~x13 & ~x15 & x10 & ~x11))))) | (x07 & ((~x15 & (x14 ? ((~x06 & (x12 | (~x10 & ~x11 & ~x12 & ~x13))) | (~x10 & ~x12 & (x11 | (x09 & ~x11 & x13)))) : (x13 ? (x10 | (~x10 & (x11 | (x09 & ~x11)))) : ~x12))) | (~x06 & ((x12 & ~x13 & (~x14 | (x14 & x15))) | (x13 & x15))) | (~x12 & ~x13 & x15))) | (x14 & ~x15 & ~x12 & ~x13 & ~x06 & ~x07 & ~x09))) | (~x04 & ~x06 & (x07 ? ~x09 : ((~x10 & (x11 | (~x09 & ~x11))) | (~x09 & x10 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))))))) | (~x05 & (x04 ? ((~x06 & ~x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))))) | (x07 & ((x12 & ((x15 & ((~x13 & x14 & (x06 ? (~x09 & (~x10 ^ ~x11)) : (x10 | (~x10 & x11)))) | (~x06 & x13 & (x10 | (~x10 & (x11 | (~x11 & (x09 | (~x09 & ~x14))))))))) | (~x06 & (x10 ? (x14 ? ~x15 : ~x13) : ((x13 & x14 & ~x09 & ~x11) | (x11 & ~x13 & ~x14)))))) | (~x06 & ((~x10 & (x11 ? ((~x12 & ~x13 & (x15 | (~x14 & ~x15))) | (~x15 & (x14 | (x13 & ~x14)))) : (x09 ? (~x15 | (~x13 & x15)) : ~x13))) | (x13 & ((~x12 & x15) | (x10 & ~x14 & ~x15))) | (x10 & ~x12 & ~x13 & (x15 | (~x14 & ~x15)))))))) : (x06 & ((~x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))))) | (~x10 & ~x11 & x07 & ~x09))))) | (x04 & x07 & ((~x09 & ((x12 & ((x06 & ~x13 & x14 & x15 & (~x10 ^ x11)) | (x13 & ~x14 & ~x15 & ~x06 & ~x10 & ~x11))) | (~x12 & x13 & ~x15 & ~x06 & ~x10 & ~x11))) | (~x12 & x14 & ~x15 & ~x06 & x10))));
  assign z17 = ~x00 & ~x01 & ~x02 & ~x03 & x09 & ((x05 & (((~x11 | (x10 & x11)) & ((x04 & x06 & x07 & x12 & x13 & x15) | (~x07 & x08 & ~x04 & ~x06))) | (x04 & ((x06 & ((~x08 & (x10 ? ((x14 & ((~x15 & (~x12 | (x12 & x13)) & (~x11 | (x07 & x11))) | (~x13 & x15 & ~x11 & x12))) | (~x13 & ~x14 & ~x11 & x12)) : ((x11 & ((~x07 & (x12 ? (x13 & ~x14) : (x14 & x15))) | (x12 & x14 & (x13 ^ x15)))) | (x07 & ~x11 & (x12 ? (x13 ? (x14 & ~x15) : ~x14) : (x14 & ~x15)))))) | (x12 & x14 & ((~x10 & x11 & x13 & x15) | (~x13 & ~x15 & x10 & ~x11))) | (x07 & ((x14 & ((~x15 & ((x10 & ((x08 & ~x12) | (x11 & x12 & ~x13))) | (~x10 & x12 & ~x13) | (x08 & ((x12 & x13) | (~x10 & ~x11 & ~x12 & ~x13))))) | (~x13 & x15 & x08 & x12))) | (~x12 & x13 & x15) | (x12 & ~x14 & ((x11 & (~x13 | (~x10 & x13 & x15))) | (x08 & ~x11 & ~x13))))))) | (x07 & ((~x06 & ((x12 & ~x13 & (~x14 | (x14 & x15))) | (x13 & x15))) | (~x12 & ~x13 & x15) | (~x15 & ((~x12 & ((~x13 & ~x14) | (~x10 & x14 & (x11 | (x08 & ~x11 & x13))))) | (x13 & ~x14) | (~x06 & x12 & x14))))) | (x14 & ~x15 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08))) | (~x04 & ~x06 & (x07 ? ~x08 : ((~x10 & (x11 | (~x08 & ~x11))) | (~x08 & x10 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))))))) | (~x05 & (x04 ? ((x07 & ((x12 & ((~x13 & ((x14 & x15 & (x06 ? (~x08 & (~x10 ^ ~x11)) : (x10 | (~x10 & x11)))) | (~x06 & ~x14 & (x10 | (~x10 & (x11 | (~x08 & ~x11 & ~x15))))))) | (~x06 & (x10 ? (x14 & ~x15) : (~x11 & (x08 ? (~x15 | (x13 & x15)) : (x14 & ~x15))))))) | (~x06 & (x10 ? ((x13 & (x15 | (~x14 & ~x15))) | (~x12 & ~x13 & x15)) : (x11 ? ((x13 & (x15 | (~x14 & ~x15))) | (x14 & ~x15) | (~x12 & ~x13 & x15)) : (x08 ? (x13 ? ~x12 : x15) : (x15 | (x13 & ~x14 & ~x15)))))))) | (~x06 & ((~x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : x15)))) | (~x14 & ~x15 & ~x12 & ~x13)))) : (x06 & ((~x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))))) | (~x10 & ~x11 & x07 & ~x08))))) | (x04 & x07 & x14 & ((~x08 & ((~x12 & x13 & ~x15 & ~x06 & ~x10 & ~x11) | (x06 & x12 & ~x13 & x15 & (~x10 ^ x11)))) | (~x06 & ~x12 & ~x15 & (x10 | (~x10 & ~x11 & ~x13))))));
  assign z18 = ~x00 & ~x01 & ~x02 & ~x03 & x10 & ((~x06 & (x04 ? ((~x15 & (x07 ? ((~x12 & ((~x09 & ((x05 & ~x08 & (x13 ? ~x11 : x14)) | (x08 & (x14 | (~x05 & ~x13 & ~x14))))) | (~x05 & (x14 | (~x13 & ~x14)) & (x11 ? ~x08 : x09)) | (x05 & x09 & x14))) | (~x14 & ((x08 & ((~x09 & x13) | (~x05 & x09 & x11 & x12))) | (~x11 & x13 & (x09 | (~x08 & ~x09 & x12))))) | (x12 & x14 & (x05 | (~x05 & (~x13 | (x13 & (~x11 | (x08 & x11)))))))) : ((~x12 & ~x13 & (x05 ? (x14 & (~x08 ^ ~x09)) : ~x14)) | (~x05 & (x14 | (x13 & ~x14)))))) | (x07 & ((x12 & ((~x13 & (x05 ? (~x14 | (x14 & x15)) : (~x14 & (~x11 | (x11 & (~x08 | (x08 & (~x09 | (x09 & x15))))))))) | (~x05 & x13 & ((x08 & x09 & x11 & x15) | (~x08 & ((x11 & x14) | (~x09 & ~x11 & x15))))))) | (~x05 & ((x15 & (((x13 | (~x12 & ~x13)) & (x09 ? ~x11 : x08)) | (~x08 & x11 & ~x12 & (~x13 | (x13 & x14))))) | (~x08 & ((~x09 & ~x11 & ~x12) | (x11 & x13 & ~x14))) | (x11 & ~x12 & x08 & x09))))) | (~x05 & ((~x13 & ((~x07 & (x12 ? ~x14 : x15)) | (x12 & x14 & x15))) | (~x07 & x13 & x15)))) : (x05 & (x07 ? (~x08 ^ ~x09) : ((x08 & x09) | ((~x08 | (x08 & ~x09)) & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))))))) | (x06 & ((x12 & ((~x13 & (((~x14 | (x14 & x15)) & (x04 ? (x05 & ((x07 & (x08 ^ ~x09)) | (~x11 & (~x08 ^ ~x09)))) : (~x05 & ~x07))) | (x04 & ((x07 & (((~x08 ^ ~x09) & ((x11 & (x14 ? x15 : x05)) | (x14 & x15 & ~x05 & ~x11))) | (x14 & ~x15 & x05 & x11))) | (x14 & ~x15 & x05 & ~x11))))) | (x04 & x05 & x13 & x14 & ~x15 & ((x07 & (x08 ^ ~x09)) | ((~x08 ^ ~x09) & (~x11 | (x07 & x11))))))) | (~x04 & ~x05 & ((~x07 & ((x14 & ~x15) | ((x15 | (~x14 & ~x15)) & (x13 | (~x12 & ~x13))))) | (x07 & ~x08 & ~x09 & ~x11))) | (x04 & x05 & ~x15 & ((x07 & ((~x12 & x14 & (x08 ? (x09 | (~x09 & x11)) : (x09 ? x11 : (~x11 | (x11 & ~x13))))) | (x13 & ~x14 & (~x11 | (x08 & ~x09 & x11))))) | (~x11 & ~x12 & x14 & (~x08 ^ ~x09)))))) | (x04 & x05 & x07 & ((~x12 & ~x13 & (x15 | (~x14 & ~x15))) | (x13 & (x15 | (x11 & ~x15 & (x08 ? (x09 & ~x14) : (~x14 | (~x09 & ~x12 & x14)))))))));
  assign z19 = ~x00 & ~x01 & ~x02 & ~x03 & x11 & ((~x06 & (x04 ? ((~x13 & ((~x12 & ((~x15 & ((~x07 & (x05 ? (x14 & (~x08 ^ ~x09)) : ~x14)) | (~x05 & x07 & ((~x08 & x10 & (~x14 | (~x09 & x14))) | (~x14 & (x09 ? ~x10 : x08)))))) | (~x05 & x15 & (~x07 | (x07 & ((x08 & (~x09 | (x09 & x10 & x14))) | (x09 & (~x10 | (~x08 & x10))) | (~x08 & ~x09 & (x14 | (x10 & ~x14))))))))) | (x07 & ((x12 & ((~x14 & ((x05 & (x09 | (~x08 & ~x09 & ~x15))) | (x08 & (~x09 | (~x05 & x09 & x10 & x15))) | (~x05 & (x10 ? ~x08 : x09)) | (~x08 & ~x09 & ~x10 & x15))) | (~x05 & ~x15 & ((x08 & (x09 ? x10 : x14)) | (~x10 & (x09 ? x14 : ~x08)))) | (x05 & x14 & x15))) | (x05 & ~x08 & ~x09 & x10 & ~x14 & x15))) | (~x05 & x12 & (x14 ? x15 : ~x07)))) | (x07 & ((x05 & ((x13 & x15) | (x12 & x14 & ~x15))) | (~x05 & ((x13 & ((~x09 & ((~x14 & (x08 ? (~x15 | (~x12 & x15)) : (x12 & ~x15))) | (~x08 & x10 & ~x12 & ~x15))) | (~x14 & (x10 ? ((x15 | (x09 & ~x15)) & (~x08 | (x08 & x12))) : ((x12 & x15) | (x09 & (~x15 | (~x12 & x15)))))) | (x14 & (x15 | (x12 & ~x15 & (~x10 | (x08 & x10))))))) | (~x08 & ((~x09 & ~x10 & ~x12 & ~x14) | (x14 & ~x15 & x10 & x12))) | (x09 & x10 & ~x12 & (x14 ? ~x15 : x08)))) | (~x12 & x14 & ~x15 & (x09 ? ~x10 : (x08 | (~x08 & ~x10)))))) | (~x05 & ~x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15)))))) : (x05 & (x07 ? (~x08 ^ ~x09) : ((x08 & x09) | ((~x08 | (x08 & ~x09)) & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))))))) | (x06 & (x04 ? (((~x08 ^ ~x09) & ((x05 & ((~x10 & ((~x07 & (x12 ? (x13 & ~x14) : (x14 & x15))) | (x12 & x14 & (x13 ^ x15)))) | (x13 & x14 & ~x15 & x07 & x10 & x12))) | (x07 & x12 & ~x13 & x14 & x15 & (x10 | (~x05 & ~x10))))) | (x05 & ((x07 & (x12 ? ((x14 & ((~x13 & ~x15) | ((x13 ^ x15) & (x08 ^ ~x09)))) | (~x13 & ~x14) | (x13 & x15 & (x10 | (~x10 & ~x14)))) : ((~x09 & x10 & ((~x14 & x15 & ~x08 & ~x13) | (x08 & x14 & ~x15))) | (x13 & x15) | (~x10 & x14 & ~x15)))) | (~x10 & x12 & x13 & x14 & x15)))) : (~x05 & ((~x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))))) | (~x09 & ~x10 & x07 & ~x08))))) | (x04 & x05 & x07 & ((x13 & ~x14 & ~x15) | (~x12 & ((x10 & ((x08 & (x09 ? (x14 & ~x15) : (~x13 & x15))) | (~x08 & x14 & (~x15 | (~x09 & ~x13 & x15))) | (x09 & ~x13 & x15))) | (~x13 & (x15 ? ~x10 : ~x14)))))));
  assign z20 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & (x07 ? (((~x08 ^ ~x09) & ((x05 & ~x06) | (~x10 & ~x11 & ~x05 & x06))) | (~x05 & x06 & ~x08 & ~x09 & (~x10 ^ ~x11))) : (x05 ? (~x06 & (x08 ? ((x09 & (~x11 | (x10 & x11))) | (~x10 & (x11 | (~x09 & ~x11))) | (~x09 & x10 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))) : ((~x10 & ~x11) | ((x10 | (~x10 & x11)) & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))))) : (x06 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))));
  assign z21 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & x05 & ~x06 & (x07 ? (~x08 ^ ~x09) : (x08 ? ((x09 & (~x11 | (x10 & x11))) | (~x10 & (x11 | (~x09 & ~x11))) | (~x09 & x10 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15))))))) : ((~x10 & ~x11) | ((x10 | (~x10 & x11)) & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))))))));
  assign z22 = ~x00 & ~x01 & ~x02 & ~x03 & x04 & ~x13 & x14 & (~x08 ^ ~x09) & ((~x05 & x06 & x07 & x12 & x15) | (x05 & ~x06 & ~x07 & ~x12 & ~x15));
  assign z23 = ~x00 & ~x02 & ((~x03 & ((x05 & ((x04 & (x01 ? (~x07 & ~x08 & x09 & x10 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))) : (x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))))))) | (x01 & ~x04 & x06 & ~x07 & ~x08 & x09 & x10 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))))) | (x01 & ~x05 & ~x07 & ~x08 & x09 & x10 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))))) | (x05 & ~x06 & ~x07 & x01 & x03 & x04));
  assign z24 = ~x00 & x01 & ~x02 & ~x03 & ~x07 & ~x11 & ~x12 & ((x04 & x05 & ~x06 & ~x08 & (x10 | (x09 & ~x10)) & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))) | (~x04 & ~x05 & x08 & ~x09 & ~x14 & ~x15 & ~x10 & ~x13));
  assign z25 = ~x00 & ~x01 & ~x02 & ~x03 & x04 & x05 & x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))) | (~x13 & (x12 ? (~x14 | (x14 & x15)) : (x15 | (~x14 & ~x15)))));
  assign z26 = ~x00 & ~x01 & ~x02 & ~x03 & x04 & x05 & x06 & ~x07 & ((x12 & x14 & ((~x10 & x11 & x13 & x15) | (~x13 & ~x15 & x10 & ~x11))) | ((~x08 ^ ~x09) & ((x14 & (x12 ? ((x13 ^ x15) & (~x10 ^ ~x11)) : (x10 ? (~x11 & ~x15) : (x11 & x15)))) | (x12 & ~x14 & (x10 ? (~x11 & ~x13) : (x11 & x13))))));
  assign z27 = x07 & x06 & x05 & ~x04 & ~x03 & ~x02 & x00 & x01;
  assign z28 = (~x00 & x01 & ~x02 & ((~x09 & ((~x07 & ((~x05 & (x03 ? (~x06 & (x08 ^ x10)) : (~x08 & x10 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))))) | (~x03 & x04 & x05 & ~x08 & x10 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))))) | (~x03 & x05 & x06 & ~x08 & x10 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15)) & (~x04 | (x04 & x07))))) | (x03 & x04 & ~x05 & (x07 | (x06 & ~x07))))) | (x00 & ~x01 & ~x03 & ~x07);
  assign z29 = (~x00 & x01 & ~x02 & ((~x10 & ((~x07 & ((~x05 & (x03 ? (~x06 & (~x08 ^ ~x09)) : (~x08 & x09 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))))) | (~x03 & x04 & x05 & ~x08 & x09 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))))) | (~x03 & x05 & x06 & ~x08 & x09 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15)) & (~x04 | (x04 & x07))))) | (x03 & x04 & x05 & (x07 | (x06 & ~x07))))) | (x00 & ~x01 & ~x03 & x07);
  assign z30 = ~x03 & (x00 ? ~x01 : (x01 & ~x02 & ((~x05 & x07) | (~x08 & ~x11 & ~x12 & (x09 ^ x10) & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15)) & (x05 ? (x04 ? (~x07 | (x06 & x07)) : x06) : ~x07)))));
  assign z31 = ~x00 & x01 & ~x02 & ~x07 & ((~x08 & ((~x05 & ((x03 & ~x06 & (x09 ^ x10)) | (~x09 & ~x10 & ~x03 & ~x04))) | (~x03 & ~x04 & x05 & x06 & ~x09 & ~x10))) | (x08 & ~x09 & ~x10 & x03 & ~x05 & ~x06));
  assign z32 = ~x00 & x01 & ~x02 & (x03 ? (x04 & ((x05 & ~x06 & ~x07) | (x06 & x07))) : (~x05 & x07));
  assign z33 = ~x03 & (x00 ? (~x01 & ~x06) : (x01 & ~x02 & ~x08 & ((~x11 & ~x12 & ~x13 & ~x14 & x15 & (x05 ? ((x06 & ((~x04 & (x10 ? ~x07 : x09)) | (x07 & ((~x09 & x10) | (x04 & x09 & ~x10))))) | (x04 & ~x07 & (x10 | (x09 & ~x10)))) : (~x07 & (x10 | (x09 & ~x10))))) | (x04 & ~x05 & ~x07 & ~x09 & ~x10))));
  assign z34 = ~x03 & (x00 ? (~x01 & x06) : (~x02 & ((x05 & ((~x13 & ((~x12 & ((x04 & ((x07 & ((~x01 & (x15 | (~x14 & ~x15))) | (x14 & ~x15 & ~x10 & ~x11 & ~x08 & x09 & x01 & x06))) | (x01 & ~x07 & ~x08 & ~x11 & x14 & ~x15 & (x10 | (x09 & ~x10))))) | (x01 & x06 & ~x08 & ~x11 & x14 & ~x15 & ((~x04 & (x10 ? ~x07 : x09)) | (x07 & ~x09 & x10))))) | (~x01 & x04 & x07 & x12 & (~x14 | (x14 & x15))))) | (~x01 & x04 & x07 & ((x14 & ~x15) | (x13 & (x15 | (~x14 & ~x15))))))) | (x01 & ~x07 & ~x08 & ((~x05 & ~x11 & ~x12 & ~x13 & x14 & ~x15 & (x10 | (x09 & ~x10))) | (~x09 & ~x10 & x04 & x06))))));
  assign z35 = ~x00 & x01 & ~x02 & ~x03 & ~x08 & ((~x11 & ~x12 & x13 & ~x14 & ~x15 & (x05 ? ((x06 & ((~x04 & (x10 ? ~x07 : x09)) | (x07 & ((~x09 & x10) | (x04 & x09 & ~x10))))) | (x04 & ~x07 & (x10 | (x09 & ~x10)))) : (~x07 & (x10 | (x09 & ~x10))))) | (~x07 & ~x09 & ~x10 & x04 & ~x05 & ~x06));
  assign z36 = x04 & (x00 ? (~x01 & ~x03) : (~x02 & ((~x03 & ((x07 & (x05 ? ((~x13 & ((~x12 & (x01 ? (x06 & ~x08 & ~x11 & (x09 ^ x10) & (~x14 ^ ~x15)) : (x15 | (~x14 & ~x15)))) | (~x01 & x12 & (~x14 | (x14 & x15))))) | (x13 & ((~x14 & ~x15 & (~x01 | (x01 & x06 & ~x08 & ~x11 & ~x12 & (x09 ^ x10)))) | (~x01 & x15))) | (~x01 & x14 & ~x15)) : x01)) | (x01 & ~x07 & ~x08 & ~x11 & ~x12 & (x10 | (x09 & ~x10)) & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))))) | (x01 & x03 & ~x06 & ~x07 & (x05 | (~x05 & (x08 ? (~x09 & ~x10) : (x09 ^ x10))))))));
  assign z37 = ~x04 & (x00 ? (~x01 & ~x03) : (x01 & ~x02 & ((~x08 & ((~x07 & ((~x05 & (x03 ? (~x06 & (x09 ^ x10)) : ((~x09 & ~x10) | (~x11 & ~x12 & (x10 | (x09 & ~x10)) & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15)))))) | (~x03 & x05 & x06 & (x10 ? (~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15))) : ~x09)))) | (~x03 & x05 & x06 & ~x11 & ~x12 & (x13 ? (~x14 & ~x15) : (~x14 ^ ~x15)) & ((x09 & ~x10) | (x07 & ~x09 & x10))))) | (~x05 & ((~x03 & x07) | (x08 & ~x09 & ~x10 & x03 & ~x06 & ~x07))))));
  assign z38 = x07 & ~x06 & x04 & x03 & ~x02 & ~x00 & x01;
  assign z39 = ~x07 & x06 & x04 & x03 & ~x02 & ~x00 & x01;
endmodule