module pla__mainpla ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53;
  assign z00 = x14 & ((~x20 & ~x21 & (x05 ? (x03 ? ((x00 & x01 & (x02 | (~x02 & ~x04 & ((~x08 & ~x09 & ~x10 & x11 & (x13 | (~x12 & ~x13 & ~x06 & ~x07))) | (x09 & ~x12 & ~x13))))) | (~x00 & ~x01 & ~x02 & x04)) : (x04 ? ((x02 & (x00 ? (x01 & x16) : (~x01 & (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))))))))) | (x00 & (~x01 | (x01 & ~x02 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) | (~x00 & x01 & ~x02 & x15)) : (x01 ? (x00 ? (~x02 | (x02 & ~x24)) : x02) : ~x02))) : (x00 ? (x03 & x04 & (x01 ^ ~x02)) : (~x03 & ~x04 & ((~x01 & ~x02 & (~x25 | (x25 & (~x24 | (~x15 & x24))))) | (x01 & x02 & ~x06 & ~x07 & ~x08 & ~x09 & x10 & ~x11 & ~x12 & ~x13)))))) | (~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & x21));
  assign z01 = x14 & ~x20 & ~x21 & ((~x01 & (x00 ? ((~x02 & x05 & (~x03 | (x03 & x04 & x22))) | (x04 & ~x05 & (~x03 | (x02 & x03)))) : (x02 ? (~x03 & x04 & x05 & (x17 | (~x17 & ((~x12 & ((~x11 & ((~x06 & ~x07 & ~x13 & ((~x08 & ~x09 & x10 & x15) | (x08 & ~x10 & ~x15))) | (x13 & ~x15 & (~x10 | (~x09 & x10))))) | (~x13 & ((x09 & ((x06 & x07 & (x08 ? (x10 | (~x10 & x11 & x18)) : x11)) | (x10 & (x15 | (x11 & ~x15))) | (~x08 & ~x10 & x11))) | (x08 & ((~x06 & ~x07 & ((~x09 & x10 & x11) | (~x10 & x15))) | (x10 & x11 & x07 & ~x09))) | (~x06 & ~x07 & ~x08 & ~x09 & ~x10 & x11 & x15 & ~x16))))) | (x13 & ((~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x10 & (x11 | (~x08 & x09 & ~x11 & x12))) | (x09 & ~x10 & (x11 | (~x11 & x12))) | (~x09 & ~x11 & x12))) | x06 | x15)) | (~x06 & ~x07 & x12 & ~x13))))) : ((~x04 & (x05 | (~x03 & ~x05 & ~x15 & x24 & x25))) | (x03 & x04 & x05))))) | (x01 & ((x04 & (x02 ? ((~x00 & x05) | (x00 & x03 & ~x05 & ~x25)) : ((~x03 & x05 & (x00 ? (x13 | (x09 & x10 & x11 & ~x12 & ~x13)) : x15)) | (~x00 & x03 & ~x05)))) | (x02 & x03 & ~x04 & x05))) | (x00 & x02 & ~x03 & x04 & x05));
  assign z02 = x14 & ((~x20 & ~x21 & (x01 ? ((~x00 & (x02 ? ((x04 & x05) | (~x03 & ~x04 & ~x05 & ~x06 & ~x07 & ~x11 & ~x12 & ~x13 & ~x08 & ~x09 & x10)) : (x03 & ~x05 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))))) | (x02 & x03 & ~x04 & x05) | (x00 & ((~x04 & ((~x12 & ~x13 & (x02 ? (~x03 & ~x05 & ((x09 & ((~x06 & ~x07 & ~x10 & (x08 ^ ~x11)) | (x08 & x10 & ~x11))) | (~x06 & ~x07 & ~x08 & x10 & ~x11))) : (x03 & x05 & (x09 | (~x09 & ~x10 & x11 & ~x06 & ~x07 & ~x08))))) | (~x02 & x03 & x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) | (x02 & ~x03 & x04 & x05 & x16)))) : (x05 ? (x02 ? (~x03 & x04 & (x00 | (~x00 & (x17 | (~x17 & (x13 ? (x06 | (~x10 & ~x15 & ((~x11 & x12 & x08 & x09) | (x11 & ~x16 & ~x08 & ~x09)))) : ((~x12 & ((x09 & ((x06 & x07 & (x08 ? x10 : x11)) | (~x06 & ~x07 & ~x10 & (x08 ? (x11 & ~x15) : ~x11)) | (x08 & x10 & ~x11 & ~x15))) | (~x06 & ~x07 & ~x08 & ~x15 & ((x10 & ~x11) | (x11 & ~x16 & ~x09 & ~x10))))) | (~x06 & ~x07 & x12)))))))) : ((x03 & (x00 ? (x04 & x22) : (~x04 | (x04 & x15)))) | (x00 & ~x03 & (~x04 | (x04 & ~x15))))) : ((x03 & ((x00 & (x04 | (~x02 & ~x04 & ~x06 & ~x07 & x08 & x11 & ~x12 & ~x13 & x09 & ~x10))) | (~x04 & x09 & ~x12 & ~x13 & ((~x00 & x08 & ((~x10 & x11 & ~x06 & ~x07) | (~x02 & x10 & ~x11))) | (~x02 & ~x06 & ~x07 & ~x08 & ~x11))))) | (~x00 & ~x02 & ~x03 & ~x04 & ~x25))))) | (~x19 & x21) | (~x04 & ((~x00 & x01 & ~x02 & ~x03) | (x00 & ~x01 & x05 & (x02 ^ x03)))));
  assign z03 = x14 & ((~x20 & ~x21 & ((x02 & ((~x03 & (x01 ? (x00 ? (x05 & (x04 ? x16 : ~x24)) : (~x04 & ~x05 & ~x12 & ~x13 & ((x09 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))) | (~x06 & ~x07 & ~x08 & ~x09 & x10 & ~x11)))) : ((x04 & x05 & (x00 | (~x00 & (x17 | (~x17 & (x13 ? (x06 | x15) : ((~x12 & ((~x06 & ((x09 & ((~x10 & x11 & x07 & x08) | (x10 & ~x11 & ~x15 & ~x07 & ~x08))) | (~x07 & (x08 ? ((~x09 & x10 & x11) | (~x10 & x15)) : (~x09 & x15 & (x10 ? ~x11 : (x11 & ~x16))))))) | (x09 & ((x06 & x07 & (x08 ? (x10 | (~x10 & x11 & x18)) : x11)) | (x15 & (x10 | (~x08 & ~x10 & x11))))) | (~x09 & x10 & x11 & x07 & x08))) | (~x06 & ~x07 & x12 & x16)))))))) | (x00 & ~x04 & ~x05 & ~x12 & ~x13 & ((x09 & ((~x06 & ~x07 & ~x10 & (x08 ^ ~x11)) | (x08 & x10 & ~x11))) | (~x06 & ~x07 & ~x08 & x10 & ~x11)))))) | (x03 & (x00 ? (x01 & (x04 ? (~x05 & ~x25) : x05)) : (~x01 & ~x04 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))))) | (~x00 & x01 & x04 & x05))) | (~x02 & ((x03 & ((x01 & (x00 ? (~x04 & x05 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ? ~x11 : (x11 & ~x15))))))) : (~x05 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))))) | (x00 & ~x01 & x04 & ~x05))) | (~x04 & ((x05 & (x00 ? ~x03 : ~x01)) | (~x00 & ~x01 & ~x03 & ~x05 & x25 & (~x24 | (~x15 & x24))))))) | (x00 & ~x01 & ~x03 & x04 & ~x05))) | (~x04 & x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))));
  assign z04 = x14 & ((~x20 & ~x21 & ((~x03 & (x04 ? (x05 & ((x02 & (x00 ? (~x01 | (x01 & x16)) : (~x01 & (x17 | (~x17 & ((~x12 & ((~x13 & (x09 ? ((x07 & ((x06 & (x08 ? x10 : x11)) | (~x10 & x11 & ~x06 & x08))) | (x10 & ~x15 & (x11 | (x08 & ~x11))) | (~x06 & ~x07 & ~x10 & (x08 ? ~x15 : ~x11))) : ((~x06 & ~x07 & ((~x15 & (x08 ? (x10 ? (x11 & ~x16) : ~x11) : (x10 ? ~x11 : (x11 & ~x16)))) | (x08 & x10 & x11 & x16))) | (x10 & x11 & x07 & x08)))) | (~x10 & x13 & ((~x11 & ~x15) | (~x06 & x07 & ~x08 & ~x09 & x11 & x16))))) | (x13 & (x06 | (~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (~x09 & ~x11 & x12) | (x11 & (x10 | (x09 & ~x10))))))) | (~x06 & ~x07 & x12 & ~x13 & x16))))))) | (x01 & ~x02 & (x00 ? ((x13 & (x15 | (x12 & ~x15))) | (x09 & x10 & x11 & ~x12 & ~x13 & x15)) : x15)))) : (x01 ? (x02 & (x00 ? (x05 & ~x24) : (~x05 & x09 & ~x12 & ~x13 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))))) : ((~x02 & ((x00 & x05) | (~x00 & ~x05 & ~x24 & x25))) | (x00 & x02 & ~x05 & ~x12 & ~x13 & ((x09 & ((~x06 & ~x07 & ~x10 & (x08 ^ ~x11)) | (x08 & x10 & ~x11))) | (~x06 & ~x07 & ~x08 & x10 & ~x11))))))) | (x03 & ((~x02 & ((~x01 & (x00 ? (~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) : (x05 & (~x04 | (x04 & ~x15))))) | (x00 & x01 & ~x04 & x05 & ~x06 & ~x07 & ~x08 & ~x09 & ~x12 & ~x13 & (x10 ? ~x11 : (x11 & x15))))) | (x01 & x02 & ((~x04 & x05) | (~x05 & ~x25 & x00 & x04))))) | (x02 & x04 & (x00 ? (~x01 & ~x05) : (x01 & x05))))) | (~x04 & ((~x00 & x01 & ~x02 & (~x03 | (x03 & x05))) | (x00 & ~x01 & x02 & ~x03 & x05))) | (~x19 & x20));
  assign z05 = x14 & ((~x20 & ~x21 & ((~x03 & (x04 ? ((x05 & (x00 ? (x01 ? (x02 ? ~x16 : (x15 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))) : (~x02 & x15)) : (x02 & (x01 | (~x01 & (x17 | (~x17 & ((~x06 & ((x16 & ((x07 & ((x12 & ~x13) | (~x08 & ~x09 & ~x10 & x11 & ~x12 & x13))) | (~x07 & x08 & ~x09 & x10 & ~x12 & ~x13))) | (~x13 & ((~x07 & ~x12 & ((x11 & ((~x08 & ~x09 & x10) | (~x15 & ((x08 & (~x10 | (~x09 & x10 & ~x16))) | (~x08 & ~x09 & ~x10 & ~x16))))) | (~x08 & ~x11 & (x09 ? ~x10 : (x10 & ~x15))))) | (x12 & ~x16))))) | (x09 & ((~x12 & ~x13 & ((x10 & ~x15 & (x11 | (x08 & ~x11))) | (x06 & x07 & (x08 ? x10 : x11)))) | (x13 & ~x15 & (x11 ? ~x10 : (x08 ? x10 : x12))))) | (x06 & (x13 | (x07 & x12 & ~x13))) | (~x09 & ((x11 & ((x08 & ((~x12 & ~x13 & x07 & x10) | (~x10 & x13 & ~x15))) | (~x08 & ~x10 & x13 & ~x15 & ~x16))) | (~x11 & x12 & x13 & ~x15))) | (x10 & x11 & x13 & ~x15))))))))) | (x00 & ~x01 & ~x02 & ~x05)) : ((x02 & (x00 ? ((~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x01 & ~x05) | (x01 & x05 & ~x24)) : (x01 & ~x05 & x09 & ~x12 & ~x13 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & ((~x08 & ~x11) | (x08 & ~x10 & x11 & ~x15))))))) | (~x00 & ~x01 & ~x02 & ~x05 & ~x24 & x25)))) | (x03 & (x00 ? (x01 ? ((~x06 & ~x07 & ~x08 & ~x02 & ~x04 & x05 & ~x09 & ~x10 & x11 & ~x12 & ~x13 & x15) | (x02 & x04 & ~x05 & x25)) : (x04 & (x02 ? ~x05 : (x05 & x22)))) : ((~x02 & ((x04 & (x01 ? ~x05 : (x05 & ~x15))) | (~x01 & ~x04 & ~x05 & x09 & ~x12 & ~x13 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))))) | (~x01 & x02 & ~x04 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13)))))) | (~x00 & ~x01 & ~x02 & ~x04 & x05))) | (~x19 & x21) | (~x04 & x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))));
  assign z06 = ~x14 | (x14 & ((~x20 & ~x21 & ((x05 & ((x04 & (x01 ? (~x03 & (x00 ? (x02 ? x16 : (~x15 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))) : (~x02 & ~x15))) : ((~x02 & (x00 ? (x03 ? x22 : ~x15) : (x03 ? ~x15 : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))) | (~x00 & x02 & ~x03 & (x17 | (~x17 & ((~x15 & (x11 ? ((~x12 & ((~x13 & ((~x06 & ~x07 & x08 & ~x09 & (~x10 | (x10 & ~x16))) | (x09 & (x10 | (~x08 & ~x10))))) | (~x08 & ~x09 & ~x10 & x13 & ~x16))) | (x13 & (x10 | (~x10 & (x09 | (x08 & ~x09)))))) : ((x09 & ((x08 & ((x10 & x13) | (~x06 & ~x07 & ~x10 & ~x12 & ~x13))) | (x12 & x13 & (~x10 | (~x08 & x10))))) | (x13 & ((~x09 & (x12 | (x10 & ~x12))) | (~x10 & ~x12)))))) | (~x13 & (x12 ? x07 : ((x07 & ((x06 & x09 & (x08 ? x10 : x11)) | (x08 & ~x09 & x10 & x11))) | (~x06 & ~x07 & ((~x08 & (x09 ? (~x10 & ~x11) : (x10 & x11))) | (x08 & ~x09 & x10 & x11 & x16)))))) | (x06 & x13)))))))) | (x03 & ~x04 & ((~x12 & ~x13 & (x00 ? (x01 & ~x02 & (x09 | (~x06 & ~x07 & ~x08 & x11 & ~x15 & ~x09 & ~x10))) : (~x01 & x02 & ((~x06 & ~x07 & ~x10 & x11 & (x08 ^ ~x09)) | (x10 & ~x11 & x08 & x09))))) | (~x02 & ((~x00 & ~x01) | (~x09 & ~x10 & x11 & x13 & x00 & x01 & ~x08))))))) | (~x05 & ((x03 & ((((x01 & x04) | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & ~x01 & ~x04)) & (~x02 | (x00 & x02))) | (~x02 & ~x04 & ~x11 & ~x12 & ~x13 & ((~x06 & ~x07 & ~x08 & ((~x00 & (x01 ? x09 : (~x09 & x10))) | (~x01 & x09))) | (x09 & x10 & ~x01 & x08))))) | (x02 & ~x03 & ~x04 & (x10 ? (~x11 & ~x12 & ~x13 & ((x00 & ((~x07 & ~x08 & x01 & ~x06) | (~x01 & x08 & x09))) | (x01 & x08 & x09))) : ((~x08 & ((x00 & ~x01 & ((~x09 & x11) | (~x11 & ~x12 & ~x13 & ~x06 & ~x07 & x09))) | (x01 & ~x06 & ~x07 & ~x12 & ~x13 & x09 & ~x11))) | (~x00 & x01 & ~x06 & ~x07 & x08 & x09 & x11 & ~x12 & ~x13 & ~x15)))))) | (~x00 & x01 & x02 & ~x03 & x04))) | (~x00 & x01 & ~x02 & ~x03 & ~x04 & x05)));
  assign z07 = x14 & ~x20 & ~x21 & (x02 ? (x03 ? (x00 ? (~x05 & ((x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & ~x01 & ~x04) | (x01 & x04 & ~x25))) : (~x01 & ~x04 & x09 & ~x12 & ~x13 & ((~x06 & ~x07 & x08 & ~x10 & x11) | (x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08 & ~x10)))))) : ((~x00 & ((~x13 & ((~x12 & ((~x06 & ~x07 & ((x09 & ((x01 & ~x04 & ~x05 & ((x08 & ~x10 & x11) | (~x08 & x10 & ~x11 & x15 & x17))) | (~x01 & x04 & x05 & ~x08 & ~x10 & ~x11 & ~x17))) | (~x01 & x04 & x05 & ~x17 & ((~x10 & (x08 | (x11 & ~x16 & ~x08 & ~x09))) | (~x09 & x10 & (x08 ? (~x11 ^ ~x16) : (x11 | (~x11 & x15)))))))) | (~x01 & x04 & x05 & ~x17 & ((~x09 & x10 & x11 & x07 & x08) | (x09 & ((x06 & x07 & (x08 ? x10 : x11)) | (x11 & (x10 ? ~x15 : ~x08)) | (x10 & (x15 | (x08 & ~x11 & ~x15))))))))) | (~x01 & x04 & x05 & x12 & ~x17 & (x06 ? x07 : (~x07 | (x07 & ~x16)))))) | (x04 & (x01 | (~x01 & x05 & (x17 | (x13 & ~x17 & (x06 | x15 | (~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (~x10 & ((x09 & (x11 | (~x11 & x12))) | (~x11 & ~x12))) | (x10 & x11) | (~x09 & ~x11 & (x12 | (x10 & ~x12))))))))))))) | (x00 & ((~x04 & ((x01 & ((x05 & ~x24) | (~x07 & ~x08 & ~x05 & ~x06 & x09 & x10 & ~x11 & ~x12 & ~x13))) | (~x05 & ((~x01 & ((~x10 & x11 & ~x08 & ~x09) | (~x11 & ~x12 & ~x13 & x08 & x09 & x10))) | (~x06 & ~x07 & ~x12 & ~x13 & ((~x08 & ~x11 & (x09 ^ x10)) | (~x10 & x11 & x08 & x09))))))) | (x01 & x04 & x05))) | (x09 & x10 & ~x11 & ~x12 & ~x13 & x01 & ~x04 & ~x05 & x08))) : (x03 ? (x04 ? (x00 ? (x01 & ~x05) : (~x01 & x05)) : ((~x12 & ~x13 & (x01 ? ((x00 & x05 & (x09 | (~x09 & ~x10 & x11 & ~x06 & ~x07 & ~x08))) | (~x00 & ~x05 & ~x06 & ~x07 & ~x08 & x09 & ~x11)) : (~x05 & ((x09 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))) | (~x00 & ~x06 & ~x07 & x10 & ~x11 & ~x08 & ~x09))))) | (~x09 & ~x10 & x11 & x13 & x05 & ~x08 & x00 & x01))) : (x00 ? (x04 & x05 & (~x01 | (x01 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : ((x01 & x04 & x05) | (~x01 & ~x04 & ~x05 & x15 & x24 & x25)))));
  assign z08 = ~x14 | (x14 & ((~x19 & (x20 | x21)) | (~x20 & ~x21 & (x02 ? ((~x00 & ((~x12 & ((~x13 & ((x10 & ((~x11 & ((~x04 & ((~x06 & ~x07 & ~x08 & ~x09) | (x08 & x09)) & (x01 ? (~x03 & ~x05) : (x03 & x05))) | (~x01 & ~x03 & x04 & x05 & ~x06 & ~x07 & ~x17 & (x08 ? (~x09 & ~x16) : ~x15)))) | (~x01 & ~x03 & x04 & x05 & ~x17 & ((x11 & ((x09 & ~x15) | (~x06 & ~x07 & ~x09 & (~x08 | (x08 & x16))))) | (x06 & x07 & x08 & x09))))) | (~x01 & x05 & ((x09 & ((~x06 & ~x07 & ((x03 & ~x04 & (x08 ? (~x10 & x11) : ~x11)) | (~x03 & x04 & ~x08 & ~x10 & ~x11 & ~x17))) | (~x03 & x04 & x11 & ~x17 & ((x06 & x07 & (~x08 | (x08 & ~x10))) | (~x08 & ~x10 & ~x15))))) | (~x06 & ~x07 & ~x08 & ~x09 & ~x10 & x11 & ((x03 & ~x04) | (~x03 & x04 & ~x15 & ~x16 & ~x17))))))) | (~x01 & ~x03 & x04 & x05 & x13 & ~x17 & ((~x09 & ((x10 & ~x11 & ~x15) | (~x08 & ~x10 & x11 & ((~x15 & ~x16) | (~x06 & x07 & x16))))) | (~x10 & ~x11 & ~x15))))) | (~x03 & x05 & ((~x04 & (x01 | (~x01 & ~x23))) | (~x01 & x04 & (x17 | (~x17 & ((x12 & ((~x06 & ~x13 & (~x07 ^ x16)) | (~x11 & x13 & ~x15 & (~x09 | (x09 & (~x10 | (~x08 & x10))))))) | (x13 & (x06 | (~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (x09 & ~x10))))))))))))))) | (x00 & ((x01 & ((x03 & x04) | (~x03 & ~x04 & ~x05 & ~x06 & ~x07 & ~x11 & ~x12 & ~x13 & ~x08 & x09 & ~x10))) | (~x03 & x04 & x05) | (~x05 & ((~x01 & ((x03 & x04) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x03 & ~x04))) | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & ~x03 & ~x04))))) | (x01 & ~x04 & ((x03 & x05) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x03 & ~x05)))) : ((x03 & ((~x01 & (x00 ? ((x04 & x05) | (~x06 & ~x07 & ~x04 & ~x05 & ~x08 & x09 & ~x11 & ~x12 & ~x13)) : ((x08 & x09 & ~x04 & ~x05 & ~x12 & ~x13 & x10 & ~x11) | (x04 & x05 & ~x15)))) | (~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x00 & ~x05 & x08 & x09 & ~x10 & x11) | (x10 & ~x11 & ~x08 & ~x09 & x00 & x01 & x05))))) | (x00 & ((~x03 & x05 & ((x04 & ~x15 & (~x01 | (x01 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) | (~x01 & ~x04 & ~x16))) | (~x01 & x04 & ~x05))) | (~x00 & ~x01 & ~x04 & x05)))) | (~x04 & ((~x00 & x01 & ~x02 & (~x03 | (x03 & x05))) | (x00 & ~x01 & x03 & x05)))));
  assign z09 = ~x14 | (x14 & ((~x20 & ~x21 & ((~x05 & ((~x04 & ((~x12 & ~x13 & ((~x06 & ~x07 & ((x09 & ((~x01 & ((x00 & ((~x02 & x03 & x08 & ~x10 & x11) | (~x08 & ~x11 & x02 & ~x03))) | (x02 & x03 & x08 & ~x10 & x11))) | (~x00 & ((x01 & x02 & ~x03 & ((~x08 & x10 & ~x11) | (x08 & ~x10 & x11 & x15))) | (~x08 & ~x11 & ~x02 & x03))))) | (~x08 & ~x09 & x10 & ~x11 & ((~x00 & ~x01 & ~x02 & x03) | (x00 & x02 & ~x03))))) | (x00 & x08 & x09 & x10 & ~x11 & ((x02 & ~x03) | (~x01 & ~x02 & x03))))) | (~x01 & ~x03 & ((~x09 & ~x10 & x11 & x00 & x02 & ~x08) | (~x00 & ~x02 & x15 & x24 & x25))))) | (x00 & x04 & (x01 ? (x03 & (~x02 | (x02 & x25))) : (x02 & ~x03))))) | (~x00 & x01 & x02 & ~x03 & x04) | (x05 & (x01 ? ((x00 & ((~x02 & (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (x04 & x15 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) | (x02 & ~x03 & x04 & x16))) | (~x00 & ~x02 & ~x03 & x04)) : ((x04 & ((~x02 & (x00 ? (x03 ? x22 : x15) : (x03 ? x15 : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))) | (~x00 & x02 & ~x03 & (x17 | (~x17 & (x13 ? (x06 | x15 | (~x08 & ~x09 & ~x10 & ~x15 & ~x16 & x11 & x12)) : (x12 ? (x06 ? x07 : ~x16) : ((x09 & ((x06 & x07 & (x08 ? x10 : x11)) | (x15 & (x10 | (~x08 & ~x10 & x11))) | (x08 & ~x15 & ((x10 & ~x11) | (~x10 & x11 & ~x06 & ~x07))))) | (~x06 & ~x07 & ((~x09 & (x08 ? ((~x10 & ~x11 & ~x15) | (x10 & x11 & x15 & ~x16)) : (x10 | (~x10 & x11 & ~x16)))) | (x08 & ~x10 & x15))))))))))) | (~x00 & x03 & ~x04 & (~x02 | (x02 & ~x08 & ((~x09 & ~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x09 ? ~x11 : (~x10 & x11)))))))))))) | (~x03 & ~x04 & x05 & (x00 ? (~x01 & x02) : (x01 & ~x02)))));
  assign z10 = x14 & ((~x20 & ~x21 & ((~x01 & (x03 ? (x04 ? ((x00 & (~x02 ^ ~x05)) | (~x00 & ~x02 & x05 & ~x15)) : (~x12 & ~x13 & ((~x06 & ~x07 & ((~x00 & ((x02 & ((~x10 & x11 & x08 & x09) | (x05 & ~x08 & (x09 ? ~x11 : (~x10 & x11))))) | (~x09 & x10 & ~x11 & ~x02 & ~x05 & ~x08))) | (~x05 & x09 & ((~x02 & (x08 ? (~x10 & x11) : ~x11)) | (x00 & x02 & x08 & ~x10 & x11))))) | (x09 & x10 & ~x11 & ~x02 & ~x05 & x08)))) : ((x05 & (x00 ? (x02 ? x04 : (x04 ? ~x15 : ~x16)) : (x04 ? ((x13 & (x02 ? (~x17 & ((~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (~x10 & ((x09 & (x11 | (~x11 & x12))) | (~x11 & ~x12))) | (x10 & x11) | (~x09 & ~x11 & (x12 | (x10 & ~x12))))) | x06 | (~x08 & ~x09 & ~x06 & x07 & ~x10 & x11 & ~x12 & x16))) : (~x12 | (~x08 & x09 & ~x10 & ~x11 & x12)))) | (x02 & (x17 | (~x13 & ~x17 & ((~x12 & ((x11 & ((x09 & ((x06 & x07 & (~x08 | (x08 & ~x10))) | (~x15 & (x10 | (~x08 & ~x10))))) | (x08 & ((~x06 & ~x07 & ~x15 & (~x10 | (~x09 & x10 & ~x16))) | (x07 & ~x09 & x10))) | (~x06 & ~x07 & ~x08 & ~x09 & ~x10 & ~x15 & ~x16))) | (x08 & ((~x11 & ((~x06 & ~x07 & ~x09 & (x10 | (~x10 & ~x15))) | (x09 & x10 & ~x15))) | (x09 & x10 & x06 & x07))) | (~x06 & ~x07 & ~x08 & x09 & ~x10 & ~x11))) | (x12 & x16 & ~x06 & x07)))))) : (~x02 | (x02 & ~x23))))) | (x00 & ~x05 & (x02 ? (~x04 & ((~x11 & ~x12 & ~x13 & x08 & x09 & x10) | (~x08 & ((~x09 & ~x10 & x11) | (~x11 & ~x12 & ~x13 & ~x06 & ~x07 & x09))))) : x04))))) | (x01 & (x05 ? (x03 ? ((x02 & (~x04 | (x00 & x04))) | (x00 & ~x02 & ~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ~x10 & x11 & (x13 | (~x06 & ~x07 & ~x12 & ~x13 & ~x15)))))) : (x00 ? (x04 & (x02 ? ~x16 : (~x15 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (x02 | (~x02 & x04 & ~x15)))) : ((x02 & ((x00 & ((x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & ~x03 & ~x04) | (x03 & x04 & ~x25))) | (~x03 & ((~x00 & (x04 | (~x04 & ~x06 & ~x07 & x08 & x09 & ~x10 & x11 & ~x12 & ~x13 & ~x15))) | (~x04 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))))) | (~x00 & ~x02 & x03 & ~x04 & ~x06 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x09)))) | (x00 & ~x05 & ((~x02 & x03 & x04) | (~x11 & ~x12 & ~x13 & ~x08 & ~x09 & x10 & x02 & ~x03 & ~x04 & ~x06 & ~x07))))) | (~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x05 & (x02 ^ x03)) | (~x00 & x01 & ~x02 & ~x03 & ~x05))));
  assign z11 = ~x14 | (x14 & ((~x20 & ~x21 & ((x02 & ((~x03 & ((~x00 & ((x17 & ((~x01 & x04 & x05) | (~x06 & ~x07 & ~x08 & x01 & ~x04 & ~x05 & x09 & x10 & ~x11 & ~x12 & ~x13 & x15))) | (~x12 & ((~x13 & ((~x06 & ~x07 & (x01 ? (~x04 & ~x05 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x04 & x05 & ~x17 & ((~x09 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x08 & ~x10) | (~x08 & ~x11 & (~x10 | (x09 & x10 & ~x15))))))) | (~x01 & x04 & x05 & ~x17 & ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (x11 & (x10 ? ~x15 : ~x08)) | (x10 & (x15 | (x08 & ~x11 & ~x15))))) | (x07 & ~x09 & (~x08 | ~x11 | (x08 & x11))))))) | (~x01 & x04 & x05 & x13 & ~x17 & ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10))))))) | (x05 & (~x04 | (~x01 & x04 & ~x17 & ((x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & (x15 | (~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))))))))))) | (x00 & (x04 ? x05 : ((x01 & ((~x07 & ~x08 & ~x05 & ~x06 & x09 & x10 & ~x11 & ~x12 & ~x13) | (x05 & x24))) | (~x05 & ((~x12 & ~x13 & ((~x06 & ~x07 & ~x08 & ~x09 & x10 & ~x11) | (x09 & ((~x06 & ~x07 & x08 & ~x10 & x11) | (~x01 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08 & ~x10))))))) | (~x09 & ~x10 & x11 & ~x01 & ~x08)))))) | (x01 & ~x04 & ~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08 & ~x10))))) | (x03 & (x01 ? (x04 ? x00 : x05) : (x00 ? (~x05 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) : (~x04 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13)))))) | (~x00 & x01 & x04))) | (x00 & ~x01 & ~x03 & x04 & ~x05) | (~x02 & ((~x01 & ((~x12 & ((~x13 & ((x09 & ((x11 & ((~x00 & ~x03 & x04 & x05 & (x10 | (~x08 & ~x10))) | (x03 & ~x04 & ~x05 & x08 & ~x10 & ~x06 & ~x07))) | (x03 & ~x04 & ~x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x00 & x03 & ~x04 & ~x05 & ~x06 & ~x07 & ~x08 & ~x09 & x10 & ~x11))) | (~x00 & ~x03 & x04 & x05 & x13))) | (x05 & ((~x00 & (~x04 | (~x08 & x09 & ~x03 & x04 & ~x10 & ~x11 & x12 & x13))) | (x00 & ~x03) | (x03 & x04))) | (~x04 & ~x05 & ~x00 & ~x03))) | (x01 & ((x05 & (x00 ? (x03 ? (~x04 & ((~x08 & ~x09 & ~x10 & x11 & (x13 | (~x12 & ~x13 & ~x06 & ~x07))) | (x09 & ~x12 & ~x13))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04))) | (~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))))) | (x00 & x03 & x04 & ~x05))))) | (~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21))));
  assign z12 = ~x14 | (x14 & ((~x20 & ~x21 & (x05 ? ((~x03 & ((x04 & (x00 ? (x01 ? (~x02 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))) : x02) : (x01 ? ~x02 : (x02 ? (x17 | (~x17 & ((~x06 & ((~x07 & ~x13 & (x12 ? x16 : (x08 ? (~x10 | (~x09 & x10 & ~x16)) : (~x09 & x15 & (x10 ? ~x11 : (x11 & ~x16)))))) | (~x09 & ~x10 & x07 & ~x08 & x11 & ~x12 & x13 & x16))) | (x13 & (x06 | x15 | (~x15 & ((~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & (~x10 | (x08 & x10 & ~x11))) | (x10 & x11) | (~x09 & ((~x11 & (x12 | (x10 & ~x12))) | (x08 & ~x10 & (x11 | (~x11 & ~x12))))))))) | (x09 & ~x12 & ~x13 & ((x11 & ((~x08 & ~x10) | (x10 & ~x15) | (x06 & x07 & (~x08 | (x08 & ~x10))))) | (x10 & (x15 | (x08 & ((~x11 & ~x15) | (x06 & x07)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (x00 & ~x02 & (~x01 | (x01 & ~x04))) | (x02 & ~x04 & (x01 | (~x00 & ~x01))))) | (~x02 & ((~x01 & ((~x00 & (~x04 | (x03 & x04))) | (x00 & x03 & x04 & ~x22))) | (x00 & x01 & x03 & ~x04 & ~x06 & ~x07 & ~x08 & ~x09 & ~x12 & ~x13 & (x10 ^ x11)))) | (x01 & x02 & x03)) : (x01 ? ((x03 & x04 & (~x00 | (x00 & x02 & x25))) | (~x00 & x02 & ~x03 & ~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : (x10 & ~x11)))) : ((x00 & (x02 ? ((x03 & x04) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x03 & ~x04)) : x04)) | (~x00 & ~x02 & ~x03 & ~x04))))) | (~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05))))));
  assign z13 = ~x14 | (x14 & ((~x20 & ~x21 & (x05 ? ((~x03 & ((x04 & (x00 ? (x01 ? (~x02 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))) : x02) : (x01 ? ~x02 : (x02 ? (x17 | (~x17 & ((~x06 & ((~x07 & ~x13 & (x12 ? x16 : (x08 ? (~x10 | (~x09 & x10 & ~x16)) : (~x09 & x15 & (x10 ? ~x11 : (x11 & ~x16)))))) | (~x09 & ~x10 & x07 & ~x08 & x11 & ~x12 & x13 & x16))) | (x13 & (x06 | x15 | (~x15 & ((~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & (~x10 | (x08 & x10 & ~x11))) | (x10 & x11) | (~x09 & ((~x11 & (x12 | (x10 & ~x12))) | (x08 & ~x10 & (x11 | (~x11 & ~x12))))))))) | (x09 & ~x12 & ~x13 & ((x11 & ((~x08 & ~x10) | (x10 & ~x15) | (x06 & x07 & (~x08 | (x08 & ~x10))))) | (x10 & (x15 | (x08 & ((~x11 & ~x15) | (x06 & x07)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (x00 & ~x02 & (~x01 | (x01 & ~x04))) | (x02 & ~x04 & (x01 | (~x00 & ~x01))))) | (~x02 & ((~x01 & ((~x00 & (~x04 | (x03 & x04))) | (x00 & x03 & x04 & ~x22))) | (x00 & x01 & x03 & ~x04 & ~x06 & ~x07 & ~x08 & ~x09 & ~x12 & ~x13 & (x10 ^ x11)))) | (x01 & x02 & x03)) : (x01 ? ((x03 & x04 & (~x00 | (x00 & x02 & x25))) | (~x00 & x02 & ~x03 & ~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : (x10 & ~x11)))) : ((x00 & (x02 ? ((x03 & x04) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x03 & ~x04)) : x04)) | (~x00 & ~x02 & ~x03 & ~x04))))) | (~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05))))));
  assign z14 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & (x05 ? ((~x03 & (x00 ? (~x02 | (x02 & x04)) : (x04 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x02 & (x04 ? x03 : ~x00)) | (~x00 & x02 & x03 & ~x04 & ((~x12 & ~x13 & ((x09 & ((~x06 & ~x07 & ~x10 & (x08 ^ ~x11)) | (x08 & x10 & ~x11))) | (~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (~x08 & ~x09 & ~x10 & x11 & x13)))) : ((~x04 & ((~x02 & ((~x00 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06))) | (x03 & x09 & ~x12 & ~x13 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))))) | (x00 & x02 & ((x09 & ~x12 & ~x13 & ((~x03 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (x08 & ~x10 & x11 & x03 & ~x06 & ~x07))) | (~x09 & ~x10 & x11 & ~x03 & ~x08))))) | (x00 & x04 & (~x03 | (x02 & x03)))))) | (x01 & ((x00 & ((~x04 & ((~x08 & ((~x06 & ~x07 & ~x12 & ~x13 & ((~x11 & ((x02 & ~x03 & ~x05 & (x10 | (x09 & ~x10))) | (~x02 & x03 & x05 & ~x09 & x10))) | (~x09 & ~x10 & x11 & ~x02 & x03 & x05))) | (~x09 & ~x10 & x11 & x13 & ~x02 & x03 & x05))) | (~x02 & x05 & (~x03 | (~x12 & ~x13 & x03 & x09))))) | (x02 & (x03 ? x04 : x05)) | (~x02 & ~x03 & x04 & x05 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) | (x05 & ((~x00 & ~x02 & ~x03 & x04) | (x02 & x03 & ~x04))) | (~x00 & (x04 ? (x02 | (~x02 & x03 & ~x05)) : (~x05 & ~x06 & ~x07 & ~x12 & ~x13 & ((x09 & (x02 ^ x03) & (x08 ? (~x10 & x11) : ~x11)) | (~x09 & x10 & ~x11 & x02 & ~x03 & ~x08))))) | (x09 & x10 & ~x11 & ~x12 & ~x13 & x02 & ~x03 & ~x04 & ~x05 & x08))) | (x00 & ~x05 & ((~x02 & x03 & x04) | (x02 & ~x03 & ~x04 & ~x06 & ~x07 & x11 & ~x12 & ~x13 & x08 & x09 & ~x10))) | (~x00 & x02 & ~x03 & ~x04 & x05)))));
  assign z15 = x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & (x05 ? ((~x03 & ((x00 & ~x02 & (~x01 | (x01 & ~x04))) | (x02 & ~x04 & (x01 | (~x00 & ~x01))) | (x04 & (x00 ? (x01 ? (~x02 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))) : x02) : (x01 ? ~x02 : (x02 ? (x17 | (~x17 & ((~x06 & (x07 ? ((~x08 & ~x09 & ~x10 & x11 & ~x12 & x13 & x16) | (x12 & ~x13 & ~x16)) : (~x13 & (x12 ? x16 : (x08 ? (~x10 | (~x09 & x10 & ~x16)) : ((~x09 & x15 & (x10 ? ~x11 : (x11 & ~x16))) | (x09 & x10 & ~x11 & ~x15))))))) | (x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x15 & ((x13 & ((~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & (~x10 | (x08 & x10 & ~x11))) | (x10 & x11) | (~x09 & ((~x11 & (x12 | (x10 & ~x12))) | (x08 & ~x10 & (x11 | (~x11 & ~x12))))))) | (x09 & x10 & ~x12 & ~x13 & (x11 | (x08 & ~x11))))) | (x06 & x13) | (~x13 & ((~x12 & ((x07 & ((x08 & ~x09 & x10 & x11) | (x09 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10 & x11))))) | (~x10 & x11 & ~x08 & x09))) | (x06 & x07 & x12)))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))))) | (x03 & (x01 ? (x02 | (x00 & ~x02 & ~x04 & ~x06 & ~x07 & ~x08 & ~x09 & ~x12 & ~x13 & (x10 ^ x11))) : ((~x00 & ((~x02 & x04) | (~x06 & ~x07 & x02 & ~x04 & ~x11 & ~x12 & ~x13 & ~x08 & x10))) | (x04 & ~x22 & x00 & ~x02)))) | (~x00 & ~x01 & ~x02 & ~x04)) : (x00 ? (~x01 & (x02 ? ((x03 & x04) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x03 & ~x04)) : x04)) : ((x01 & (x04 ? x03 : (~x06 & ~x07 & ~x12 & ~x13 & ((x02 & ~x03 & ((~x08 & x10 & ~x11) | (~x10 & x11 & x08 & x09))) | (x09 & ~x10 & x11 & ~x02 & x03 & x08))))) | (~x01 & ~x02 & ~x03 & ~x04))))));
  assign z16 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & ((x05 & ((~x01 & ((~x03 & (x00 ? (~x02 | (x02 & x04)) : (x04 & (x02 ? (x17 | (~x17 & ((~x06 & (x07 ? (x16 & ((x12 & ~x13) | (~x08 & ~x09 & ~x10 & x11 & ~x12 & x13))) : (~x13 & (x12 | (~x12 & (x08 ? (~x10 | (~x09 & x10)) : ((~x11 & (x09 ? (~x10 | (x10 & ~x15)) : (x10 & x15))) | (~x09 & x11 & (x10 | (~x10 & ~x16)))))))))) | (x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (x11 & ((~x12 & ~x13 & ((x06 & x07 & (x08 ? (x09 ^ x10) : x09)) | (x09 & (x10 ? ~x15 : ~x08)))) | (x13 & ~x15 & (x10 | (~x10 & (x09 | (~x09 & (x08 | (~x08 & ~x16))))))))) | (x06 & (x13 | (x07 & ~x13 & (x12 | (x08 & x09 & x10 & ~x12))))) | (~x11 & ~x15 & ((x13 & ((~x09 & (x12 | (x10 & ~x12))) | (~x10 & ~x12))) | (x09 & (x10 ? (x08 ? (x13 | (~x12 & ~x13)) : (x12 & x13)) : (x12 & x13)))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x02 & (x04 ? x03 : ~x00)) | (~x00 & x02 & x03 & ~x04 & ((~x08 & ~x09 & ~x10 & x11 & x13) | (~x12 & ~x13 & ((x09 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))) | (~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))))))) | (~x03 & (x00 ? (x01 & (x02 | (~x02 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))))) : ((x02 & ~x04) | (x01 & ~x02 & x04)))) | (x01 & x03 & ((x02 & (~x04 | (x00 & x04))) | (x00 & ~x02 & ~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))))))) | (~x05 & (x04 ? ((x03 & ((x01 & (x00 ? (x02 & ~x25) : ~x02)) | (x00 & (~x02 | (~x01 & x02))))) | (x00 & ~x01 & ~x03)) : ((~x12 & ~x13 & ((~x11 & ((x10 & ((x02 & ~x03 & ((x00 & ((~x07 & ~x08 & x01 & ~x06) | (~x01 & x08 & x09))) | (x01 & ((x08 & x09) | (~x00 & ~x06 & ~x07 & ~x08 & ~x09))))) | (~x01 & ~x02 & x03 & ((x08 & x09) | (~x00 & ~x06 & ~x07 & ~x08 & ~x09))))) | (~x06 & ~x07 & ~x08 & x09 & (x02 ? (~x03 & (x00 ? (~x01 | (x01 & ~x10)) : x01)) : (x03 & (~x01 | (~x00 & x01))))))) | (~x06 & ~x07 & x08 & x09 & ~x10 & x11 & (x02 ? (x00 ? (~x03 | (~x01 & x03)) : (x01 & ~x03)) : (x03 & (~x01 | (~x00 & x01))))))) | (~x01 & ~x03 & ((~x00 & ~x02) | (~x09 & ~x10 & x11 & x00 & x02 & ~x08)))))) | (~x00 & x01 & x02 & x04))));
  assign z17 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & (x05 ? ((~x03 & ((x00 & ~x02 & (~x01 | (x01 & ~x04))) | (x02 & ~x04 & (x01 | (~x00 & ~x01))) | (x04 & (x00 ? (x01 ? (~x02 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))) : x02) : (x01 ? ~x02 : (x02 ? (x17 | (~x17 & ((x13 & (x06 | x15 | (~x15 & ((~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & (~x10 | (x08 & x10 & ~x11))) | (x10 & x11) | (~x09 & ((~x11 & (x12 | (x10 & ~x12))) | (x08 & ~x10 & (x11 | (~x11 & ~x12))))))))) | (x09 & ~x12 & ~x13 & ((x11 & ((~x08 & ~x10) | (x10 & ~x15) | (x06 & x07 & (~x08 | (x08 & ~x10))))) | (x10 & (x15 | (x08 & ((~x11 & ~x15) | (x06 & x07))))))) | (~x06 & ((~x09 & ~x10 & x07 & ~x08 & x11 & ~x12 & x13 & x16) | (~x13 & (x07 ? ((x12 & ~x16) | (x08 & ~x09 & x10 & x11 & ~x12)) : (x12 ? x16 : (x08 ? (~x10 | (~x09 & x10 & ~x16)) : (~x09 & ((~x10 & x11 & x15 & ~x16) | (x10 & (x11 | (~x11 & x15)))))))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))))) | (~x00 & ~x01 & ~x02 & ~x04) | (x03 & (x01 ? (x02 | (x00 & ~x02 & ~x04 & ~x06 & ~x07 & ~x08 & ~x09 & ~x12 & ~x13 & (x10 ^ x11))) : ((x04 & ~x22 & x00 & ~x02) | (~x00 & ((~x02 & x04) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & x02 & ~x04))))))) : ((~x01 & ((x00 & (x02 ? ((x03 & x04) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x03 & ~x04)) : x04)) | (~x00 & ~x02 & ~x03 & ~x04))) | (~x00 & x01 & ((x03 & x04) | (x02 & ~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x08 & x10 & ~x11) | (~x10 & x11 & x08 & x09)))))))));
  assign z18 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & (x05 ? ((~x03 & ((~x04 & (x00 ? (x01 & ~x02) : x02)) | (x04 & (x00 ? (x01 ? (~x02 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))) : x02) : (x01 ? ~x02 : (x02 ? (x17 | (~x17 & ((x13 & (x06 | x15 | (~x15 & ((~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & (~x10 | (x08 & x10 & ~x11))) | (x10 & x11) | (~x09 & ((~x11 & (x12 | (x10 & ~x12))) | (x08 & ~x10 & (x11 | (~x11 & ~x12))))))))) | (x09 & ~x12 & ~x13 & ((x11 & ((~x08 & ~x10) | (x10 & ~x15) | (x06 & x07 & (~x08 | (x08 & ~x10))))) | (x10 & (x15 | (x08 & ((~x11 & ~x15) | (x06 & x07))))))) | (~x06 & (x07 ? (x16 & ((x12 & ~x13) | (~x08 & ~x09 & ~x10 & x11 & ~x12 & x13))) : (~x13 & (x12 | (~x12 & ((x08 & ~x10) | (~x09 & ((~x08 & ~x10 & x11 & ~x16) | (x10 & (x08 ? (x11 | (~x11 & ~x16)) : (~x11 & x15)))))))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (x00 & (x01 ^ ~x02)))) | (x03 & (x04 ? ((~x01 & ~x02) | (x00 & x01 & x02)) : ((~x12 & ~x13 & ((~x06 & ~x07 & ~x08 & ((x00 & x01 & ~x02 & ~x09 & (x10 ^ x11)) | (x09 & ~x10 & ~x11 & ~x00 & ~x01 & x02))) | (x10 & ~x11 & x08 & x09 & ~x00 & ~x01 & x02))) | (x01 & (x02 | (~x09 & ~x10 & x11 & x13 & x00 & ~x02 & ~x08)))))) | (~x00 & (x01 ? (x02 & x04) : (~x02 & ~x04)))) : ((x04 & (x00 ? ~x01 : (x01 & x03))) | (~x03 & ~x04 & ((~x00 & ~x01 & ~x02) | (x02 & ~x12 & ~x13 & ((~x06 & ~x07 & (x00 ? (~x01 & ((~x08 & x10 & ~x11) | (~x10 & x11 & x08 & x09))) : (x01 & ((~x10 & x11 & x08 & x09) | (~x08 & ~x11 & (x09 | (~x09 & x10))))))) | (x09 & x10 & ~x11 & x00 & x01 & x08)))))))));
  assign z19 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & ((x05 & ((~x01 & ((~x03 & (x00 ? (~x02 | (x02 & x04)) : (x04 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x10 & ((~x12 & ((x11 & ((~x08 & ((~x06 & ~x09 & (x07 ? (x13 & x16) : (~x13 & ~x16))) | (x09 & ~x13))) | (x06 & x07 & x08 & x09 & ~x13))) | (~x06 & ~x07 & ~x13 & (x08 | (~x08 & x09 & ~x11))) | (x08 & ~x09 & ~x11 & x13 & ~x15))) | (x13 & ~x15 & (x09 | (~x09 & x11 & (x08 | (~x08 & ~x16))))))) | (x10 & ((~x12 & ((~x13 & ((~x06 & ~x07 & (~x09 | (~x11 & ~x15 & ~x08 & x09))) | (x08 & ((x09 & ~x11 & ~x15) | (x07 & (x09 ? x06 : x11)))) | (x09 & x11 & ~x15))) | (x13 & ~x15 & ~x09 & ~x11))) | (x13 & ~x15 & (x11 | (x09 & ~x11 & (x08 | (~x08 & x12))))))) | (x06 & (x13 | (x07 & ~x13 & (x12 | (~x08 & x09 & x11 & ~x12))))) | (x12 & ((x13 & ~x15 & ~x09 & ~x11) | (~x06 & ~x13)))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x02 & (x04 ? x03 : ~x00)) | (~x00 & x02 & x03 & ~x04 & ~x08 & ((~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))) | (~x06 & ~x07 & x09 & ~x12 & ~x13 & ~x10 & ~x11))))) | (~x03 & (x00 ? (x01 & (x02 | (~x02 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))))) : ((x02 & ~x04) | (x01 & ~x02 & x04)))) | (x01 & x03 & (x02 | (x00 & ~x02 & ~x04 & ~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))))) | (~x05 & (x04 ? ((x01 & ((~x00 & (x02 | (~x02 & x03))) | (x00 & x02 & x03 & ~x25))) | (x00 & ((~x02 & x03) | (~x01 & (~x03 | (x02 & x03)))))) : ((~x01 & ~x03 & ((~x00 & ~x02) | (~x09 & ~x10 & x11 & x00 & x02 & ~x08))) | (~x06 & ~x07 & ~x12 & ~x13 & ((x09 & (x00 ? ((~x01 & ((~x10 & x11 & x03 & x08) | (~x08 & x10 & ~x11 & x02 & ~x03))) | (x02 & ~x03 & x08 & ~x10 & x11)) : ((~x08 & ~x11 & ~x02 & x03) | (x01 & ((~x02 & x03 & x08 & ~x10 & x11) | (x02 & ~x03 & (x08 ? (~x10 & x11) : ~x11))))))) | (~x08 & ~x09 & x10 & ~x11 & (x00 ? (x02 & ~x03) : (x01 ? (x02 & ~x03) : (~x02 & x03))))))))) | (x03 & ~x04 & ~x06 & ~x00 & ~x01 & x02 & ~x07 & x08 & x09 & ~x12 & ~x13 & ~x10 & x11))));
  assign z20 = x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & (x05 ? ((~x03 & (x00 ? (x01 & (x02 | (~x02 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))))) : ((x02 & ~x04) | (x01 & ~x02 & x04)))) | (x01 & x03 & (x02 | (x00 & ~x02 & ~x04 & ~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) | (~x01 & ((~x03 & (x00 ? (~x02 | (x02 & x04)) : (x04 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & ((~x13 & ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10 & x11))) | (x10 & ~x15 & (x11 | (x08 & ~x11))) | (~x08 & ~x10 & x11))) | (~x09 & x10 & x11 & x07 & x08) | (~x06 & ~x07 & ((x08 & ~x10) | (~x09 & ((~x08 & ~x10 & x11 & ~x16) | (x10 & (~x08 | (x08 & (x11 | (~x11 & ~x16))))))))))) | (~x09 & x13 & (x10 ? (~x11 & ~x15) : ((x08 & ~x11 & ~x15) | (~x06 & x07 & ~x08 & x11 & x16)))))) | (x06 & (x13 | (x07 & x12 & ~x13))) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & ~x10) | (x10 & x11) | (~x09 & ~x11 & x12))) | (~x06 & x12 & ~x13)))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x02 & (x04 ? x03 : ~x00)) | (~x00 & x02 & x03 & ~x04 & ~x08 & ((~x11 & ~x12 & ~x13 & ~x06 & ~x07 & x09) | (~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11))))))))) : ((x02 & (x00 ? (x03 ? (x01 ? (x04 & ~x25) : (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) : (~x04 & ((~x08 & ((~x01 & ((~x09 & ~x10 & x11) | (~x06 & ~x07 & x09 & ~x12 & ~x13 & x10 & ~x11))) | (~x12 & ~x13 & x10 & ~x11 & ~x06 & ~x07 & ~x09))) | (~x12 & ~x13 & ~x10 & x11 & ~x06 & ~x07 & x08 & x09)))) : (x01 & (x04 | (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (~x08 & ~x11 & (x09 | (~x09 & x10))))))))) | (x04 & ((~x00 & x01 & ~x02 & x03) | (x00 & (x03 ? ~x02 : ~x01)))) | (~x00 & ~x02 & ~x04 & (x01 ? (x03 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)) : ~x03))))));
  assign z21 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & (x05 ? ((~x03 & (x01 ? (x02 ? (~x04 | (x00 & x04 & x16)) : (x00 ? (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))) : x04)) : (x00 ? (~x02 | (x02 & x04)) : (x04 ? (x02 ? (x17 | (~x17 & ((~x06 & ((x07 & ((~x08 & ~x09 & ~x10 & x11 & ~x12 & x13 & x16) | (x12 & ~x13 & ~x16))) | (~x13 & ((x12 & x16) | (~x07 & ~x12 & (x08 ? (~x10 | (~x09 & x10)) : (x09 ? (~x10 & ~x11) : ((~x10 & x11 & x15 & ~x16) | (x10 & (x11 | (~x11 & x15))))))))))) | (x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x15 & ((x13 & ((~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & (~x10 | (x08 & x10 & ~x11))) | (x10 & x11) | (~x09 & ((~x11 & (x12 | (x10 & ~x12))) | (x08 & ~x10 & (x11 | (~x11 & ~x12))))))) | (x09 & x10 & ~x12 & ~x13 & (x11 | (x08 & ~x11))))) | (x06 & x13) | (~x13 & ((x06 & x07 & x12) | (~x12 & ((~x09 & x10 & x11 & x07 & x08) | (x09 & ((~x08 & ~x10 & x11) | (x06 & x07 & (x08 ? (x10 | (~x10 & x11)) : x11))))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))) : x02)))) | (~x00 & ~x01 & ~x02 & ~x04) | (x03 & (x01 ? (x02 | (x00 & ~x02 & ~x04 & ~x06 & ~x07 & ~x08 & ~x09 & ~x12 & ~x13 & (x10 ^ x11))) : ((x04 & ~x22 & x00 & ~x02) | (~x00 & ((~x02 & x04) | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & x02 & ~x04))))))) : (x04 ? ((x03 & (x00 ? (x02 & (~x01 | (x01 & ~x25))) : x01)) | (x00 & ~x01 & ~x02)) : ((~x06 & ~x07 & ~x12 & ~x13 & ((x09 & ((~x01 & ((x00 & ((~x02 & x03 & x08 & ~x10 & x11) | (~x08 & x10 & ~x11 & x02 & ~x03))) | (~x08 & ~x10 & ~x11 & ~x00 & ~x02 & x03))) | (~x00 & x01 & x02 & ~x10 & x11 & ~x03 & x08))) | (~x00 & x01 & x02 & x10 & ~x11 & ~x03 & ~x08))) | (~x00 & ~x01 & ~x02 & ~x03))))));
  assign z22 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & ((~x03 & ((x05 & (x01 ? (x02 ? (~x04 | (x00 & x04 & x16)) : (x00 ? (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))) : x04)) : (x00 ? (~x02 | (x02 & x04)) : (x04 ? (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x15 & ((x13 & ((~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & (~x10 | (x08 & x10 & ~x11))) | (x10 & x11) | (~x09 & ((~x11 & (x12 | (x10 & ~x12))) | (x08 & ~x10 & (x11 | (~x11 & ~x12))))))) | (x09 & x10 & ~x12 & ~x13 & (x11 | (x08 & ~x11))))) | (x06 & x13) | (~x13 & ((x06 & x07 & x12) | (~x12 & ((~x09 & x10 & x11 & x07 & x08) | (x09 & ((~x08 & ~x10 & x11) | (x06 & x07 & (x08 ? (x10 | (~x10 & x11)) : x11)))))))) | (~x06 & ((x07 & ((~x08 & ~x09 & ~x10 & x11 & ~x12 & x13 & x16) | (x12 & ~x13 & ~x16))) | (~x13 & ((x12 & x16) | (~x07 & ~x12 & (x08 ? (~x10 | (~x09 & x10)) : ((x09 & x10 & ~x11 & ~x15) | (~x09 & ((~x10 & x11 & x15 & ~x16) | (x10 & (x11 | (~x11 & x15))))))))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))) : x02)))) | (~x04 & ~x05 & ((~x00 & ~x01 & ~x02) | (x02 & ~x12 & ~x13 & ((~x06 & ~x07 & ((~x08 & ~x11 & ((x09 & ((x00 & (~x01 | (x01 & ~x10))) | (x01 & x10))) | (~x09 & x10 & ~x00 & x01))) | (x09 & ~x10 & x11 & ~x00 & x01 & x08))) | (x09 & x10 & ~x11 & x00 & ~x01 & x08))))))) | (x03 & ((~x02 & ((~x04 & ~x12 & ~x13 & ((~x06 & ~x07 & ~x08 & ((x00 & x01 & x05 & ~x09 & (x10 ^ x11)) | (~x00 & ~x01 & ~x05 & x10 & ~x11))) | (x10 & ~x11 & x08 & x09 & ~x00 & ~x01 & ~x05))) | (~x01 & x04 & x05 & (~x00 | (x00 & ~x22))))) | (x02 & ((x01 & x05) | (x00 & x04 & ~x05 & (~x01 | (x01 & ~x25))))) | (~x00 & x01 & x04 & ~x05))) | (~x01 & ~x02 & (x00 ? (x04 & ~x05) : (~x04 & x05))))));
  assign z23 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x00 & ((~x01 & ((~x04 & (x02 ? (x03 & ((x05 & ~x08 & ~x09 & ~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & ((x09 & ((x08 & ~x10 & x11) | (x05 & ~x08 & ~x11))) | (x05 & ~x08 & ~x09 & (x10 ^ x11)))))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x09 & (x10 ? (~x11 & ~x15) : ((x08 & ~x11 & ~x15) | (x07 & ~x08 & x11 & (~x16 | (~x06 & x16)))))) | (x10 & ~x11 & ~x08 & x09)) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15))) | (~x09 & ~x10 & x07 & ~x08)) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x10 & x11) | (~x10 & (x09 | (x11 & ~x16 & ~x08 & ~x09)))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x03 & ((x05 & ((x02 & ~x04) | (x01 & ~x02 & x04))) | (x01 & x02 & ~x04 & ~x05 & ~x12 & ~x13 & ((x09 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))) | (~x06 & ~x07 & ~x08 & ~x09 & x10 & ~x11))))) | (x01 & (x02 ? x04 : (x03 & ~x05 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))))) | (~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x09 & ~x02 & x03 & ~x04 & ~x05 & ~x06))) | (x00 & ((~x02 & ((~x01 & ((~x03 & x05) | (x09 & x10 & ~x11 & ~x12 & ~x13 & ~x05 & x08 & x03 & ~x04))) | (x01 & x05 & (x03 ? (~x04 & ~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))))) | (x03 & x04 & ~x05))) | (x02 & ((x01 & (x03 ? x04 : x05)) | (~x01 & ((x04 & (~x03 ^ ~x05)) | (~x03 & ~x04 & ~x05 & ~x08 & ((~x09 & ~x10 & x11) | (~x06 & ~x07 & x09 & ~x12 & ~x13 & x10 & ~x11))))) | (~x03 & ~x04 & ~x05 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))))) | (~x01 & ~x05 & ((~x03 & x04) | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & x03 & ~x04))))) | (x03 & x05 & (x01 ? (x02 & ~x04) : (~x02 & x04)))))));
  assign z24 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & ((~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))) | (x12 & ((~x06 & ~x13) | (x07 & (x13 ? ((~x08 & (x09 ? (x10 & ~x11) : ~x10)) | (x10 & ~x11 & x08 & ~x09)) : x06))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))))) | (x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04)))))));
  assign z25 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x07 & (x09 ? ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11)) : (~x08 | ~x11 | (x08 & x11)))) | (x08 & ((~x06 & ~x07 & ~x10) | (x09 & x10 & ~x11 & ~x15))) | (~x08 & ((x09 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (~x06 & ~x07 & ~x10 & (~x11 | (~x09 & x11 & ~x16))))) | (~x06 & ~x07 & ~x09 & x10)))) | (x12 & (x13 ? ((~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15))) | (~x09 & ~x10 & x07 & ~x08)) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (~x08 & ~x09 & ~x10 & x11 & x13 & ~x15 & ~x16)))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z26 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & ((~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((~x12 & ((~x13 & ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (x10 & (x15 | (x11 & ~x15))) | (~x08 & ((~x06 & ~x07 & x10 & ~x11 & ~x15) | (~x10 & x11 & x15))))) | (~x09 & ((x07 & (~x08 | ~x11 | (x08 & ~x10 & x11))) | (~x06 & ~x07 & (x08 ? ((x11 & (x10 ? (x15 & ~x16) : ~x15)) | (x10 & (x16 | (~x11 & ~x16)))) : (x10 ? (x11 | (~x11 & x15)) : (~x11 | (x11 & x15 & ~x16))))))) | (~x06 & ~x07 & x08 & ~x10 & x15))) | (~x08 & x13 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & (x15 | (~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (x09 & ~x10)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (((~x02 & x03) | (x00 & x02 & ~x03)) & ((x04 & x05) | (x08 & x09 & ~x04 & ~x05 & ~x12 & ~x13 & x10 & ~x11))) | (x00 & ((~x02 & ((~x03 & x05) | (~x11 & ~x12 & ~x13 & ~x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (~x05 & ((~x03 & x04) | (x02 & (x03 ? (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06)) : (~x04 & ~x08 & ((~x09 & ~x10 & x11) | (~x11 & ~x12 & ~x13 & ~x06 & ~x07 & x09))))))))) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & ~x02 & x03 & ~x04))) | (x01 & ((x00 & (x02 ? (x03 ? (x04 & (x05 | (~x05 & x25))) : (x05 | (~x06 & ~x07 & ~x08 & ~x04 & ~x05 & ~x11 & ~x12 & ~x13 & x09 & ~x10))) : (x05 & (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))))))) | (x05 & ((~x00 & ~x02 & ~x03 & x04) | (x02 & x03 & ~x04))) | (~x05 & (x02 ? (~x03 & ~x04 & ~x12 & ~x13 & ((~x00 & ~x06 & ~x07 & x10 & ~x11 & ~x08 & ~x09) | (x09 & ((x08 & x10 & ~x11) | (~x00 & ~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))))) : (x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & ~x00 & ~x04))))) | (~x00 & x02 & x04))) | (~x04 & ((x02 & ~x03 & (x00 ? (~x05 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : x05)) | (~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x09 & ~x00 & ~x02 & x03 & ~x05 & ~x06)))))));
  assign z27 = x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((x02 & ((~x03 & ((~x00 & ((x05 & (~x04 | (~x01 & x04 & (x17 | (~x17 & ((~x06 & ((~x09 & ~x10 & x07 & ~x08 & x11 & ~x12 & x13 & x16) | (~x13 & ((x07 & ((x12 & ~x16) | (x08 & x09 & ~x10 & x11 & ~x12))) | (x12 & x16) | (~x07 & ~x12 & (x10 ? ~x09 : (x08 ? (x15 | (~x15 & (x09 | (~x09 & ~x11)))) : (~x11 | (~x09 & x11 & ~x16))))))))) | (x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (x13 & ((~x09 & ((x08 & ((~x10 & x11 & ~x15) | (~x11 & x12 & x07 & x10))) | (~x08 & ~x10 & ((x07 & (x12 | (x11 & ~x12 & ~x16))) | (x11 & ~x15 & ~x16))) | (~x11 & ~x15 & (x12 | (x10 & ~x12))))) | (~x15 & (x11 ? (x10 | (x09 & ~x10)) : ((~x10 & ~x12) | (x09 & (x10 ? (x08 | (~x08 & x12)) : x12))))) | x06 | (~x08 & x09 & x10 & ~x11 & (~x12 | (x07 & x12))))) | (~x13 & ((x06 & x07 & x12) | (~x12 & ((x07 & ~x09 & (~x08 | ~x11 | (x08 & x11))) | (x09 & ((x10 & ((x11 & ~x15) | (x08 & ((~x11 & ~x15) | (x06 & x07))))) | (~x08 & ~x10 & x11) | (x07 & ((x06 & x11 & (~x08 | (x08 & ~x10 & ~x18))) | (~x11 & (~x08 | (x08 & ~x10))))))))))) | (x06 & ~x07))))))) | (x01 & ~x04 & ~x05 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (~x08 & ~x11 & (x09 | (~x09 & x10))))))) | (~x04 & ((x00 & ((x01 & ((~x07 & ~x08 & ~x05 & ~x06 & x09 & x10 & ~x11 & ~x12 & ~x13) | (x05 & x24))) | (~x05 & ((~x09 & ~x10 & x11 & ~x01 & ~x08) | (~x12 & ~x13 & ((~x11 & ((~x01 & x10 & ((~x06 & ~x07 & ~x08) | (x08 & x09))) | (~x06 & ~x07 & ~x08 & x09 & ~x10))) | (~x06 & ~x07 & x08 & x09 & ~x10 & x11))))))) | (~x12 & ~x13 & x10 & ~x11 & x08 & x09 & x01 & ~x05))))) | (x03 & (x01 ? ((~x04 & x05) | (~x05 & ~x25 & x00 & x04)) : (x00 ? (~x05 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) : (~x04 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13)))))) | (x01 & x04 & (~x00 | (x00 & x05))))) | (~x02 & (x03 ? (x04 ? (x00 ? (~x05 | (~x01 & x05 & ~x22)) : (~x01 ^ ~x05)) : ((~x09 & ~x10 & x11 & x13 & x05 & ~x08 & x00 & x01) | (~x12 & ~x13 & ((~x06 & ~x07 & ((~x08 & (x01 ? ((x00 & x05 & ~x09 & (x10 ^ x11)) | (~x00 & ~x05 & x09 & ~x11)) : (~x05 & ~x11 & (x09 | (~x00 & ~x09 & x10))))) | (~x05 & x08 & x09 & ~x10 & x11 & (~x01 | (~x00 & x01))))) | (x09 & ((x00 & x01 & x05) | (x08 & x10 & ~x11 & ~x01 & ~x05))))))) : (x05 & (x04 ? ((x01 & (~x00 | (x00 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) | (~x00 & ~x01 & ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))) : (~x01 | (x00 & x01)))))) | (x00 & ~x01 & ~x03 & x04))));
  assign z28 = x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((x05 & ((~x00 & ((~x01 & (x02 ? (x03 ? (~x04 & ((~x08 & ~x09 & ~x10 & x11 & x13) | (~x12 & ~x13 & ((~x09 & ~x10 & x11 & ~x06 & ~x07 & ~x08) | (~x11 & ((x08 & x09 & x10) | (~x06 & ~x07 & ~x08 & (x09 | (~x09 & x10))))))))) : (x04 & (x17 | (~x17 & ((~x12 & ((~x09 & ((~x08 & ((~x06 & ((~x07 & ~x13 & (x10 ? (x11 | (~x11 & x15)) : (~x11 | (x11 & x15 & ~x16)))) | (x07 & ~x10 & x11 & x13 & x16))) | (x07 & (~x13 | (~x10 & x11 & x13 & ~x16))))) | (~x13 & ((x07 & (~x11 | (x08 & ~x10 & x11))) | (~x06 & ~x07 & x08 & x10 & (x16 | (~x16 & (~x11 | (x11 & x15))))))))) | (~x13 & ((x08 & ((x07 & x09 & ((x06 & (x10 | (~x10 & x11 & ~x18))) | (~x10 & (~x11 | (~x06 & x11))))) | (~x06 & ~x07 & ~x10 & x15))) | (x09 & ((x10 & x15) | (~x08 & ((~x10 & x11 & x15) | (x07 & (~x11 | (x06 & x11))))))))) | (~x08 & x09 & x10 & ~x11 & x13))) | (x12 & ((~x13 & (x06 ? x07 : (x16 | (x07 & ~x16)))) | (x07 & x13 & ((~x08 & (x09 ? (x10 & ~x11) : ~x10)) | (x10 & ~x11 & x08 & ~x09))))) | (x06 & (~x07 | x13)) | (x13 & x15)))))) : (x04 & (x03 | (~x03 & ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))) | (~x03 & ((x02 & ~x04) | (x01 & ~x02 & x04))))) | (~x02 & ((~x01 & ((~x03 & ~x04) | (x00 & x03 & x04 & ~x22))) | (x00 & x01 & (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))))))) | (x01 & x02 & ((x03 & ~x04) | (x00 & (x04 | (~x03 & ~x04 & x24))))))) | (~x05 & ((x03 & ((~x02 & ((x01 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & ~x00 & ~x04))) | (~x04 & ~x12 & ~x13 & ((~x06 & ~x07 & ((~x08 & ~x11 & ((~x00 & (x09 | (~x01 & ~x09 & x10))) | (x09 & ~x10 & x00 & ~x01))) | (~x01 & x08 & x09 & ~x10 & x11))) | (x09 & x10 & ~x11 & ~x01 & x08))))) | (x00 & ~x01 & x02 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))))) | (x02 & ~x03 & ~x04 & (x08 ? (x09 & ~x12 & ~x13 & ((x00 & ((~x10 & x11 & ~x06 & ~x07) | (~x01 & x10 & ~x11))) | (x01 & ((x10 & ~x11) | (~x00 & ~x06 & ~x07 & ~x10 & x11))))) : ((~x06 & ~x07 & ~x11 & ~x12 & ~x13 & (x00 ? (x10 ? ~x01 : x09) : (x01 & (x09 | (~x09 & x10))))) | (~x09 & ~x10 & x11 & x00 & ~x01)))))) | (x00 & ~x01 & ~x03 & x04) | (~x00 & x02 & ((x01 & x04) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x04 & ~x06 & ~x07 & ~x01 & x03))))));
  assign z29 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x06 & (~x07 | (x07 & x12 & ~x13))) | (~x12 & (x13 ? ((~x11 & ~x15 & (~x10 | (~x09 & x10))) | (~x08 & (x09 ? (x10 & ~x11) : (~x10 & x11 & ((~x15 & ~x16) | (x07 & (~x16 | (~x06 & x16)))))))) : (((x15 | (x11 & ~x15)) & ((x09 & x10) | (x08 & ~x10 & ~x06 & ~x07))) | (~x08 & ((x07 & (~x09 | (x09 & ~x11))) | (x09 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (~x06 & ~x07 & ((~x10 & ~x11) | (~x09 & (x10 ? ~x11 : (x11 & ~x16))))))) | (x08 & ((~x06 & ~x07 & ((~x09 & x10) | (~x11 & ~x15 & x09 & ~x10))) | (x09 & x10 & ~x11 & ~x15) | (x07 & (x09 ? ~x10 : x11)))) | (x07 & ~x09 & ~x11)))) | (~x06 & x12 & ~x13) | (x13 & (x15 | (~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (x09 & ~x10))))) | (x12 & ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z30 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & ((x05 & ((~x03 & (x00 ? (x01 & (x02 | (~x02 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))))) : ((x02 & ~x04) | (x01 & ~x02 & x04)))) | (x01 & x03 & ((x02 & (~x04 | (x00 & x04))) | (x00 & ~x02 & ~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))))) | (~x01 & ((~x03 & (x00 ? (~x02 | (x02 & x04)) : (x04 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))) | (~x12 & ((~x08 & ((x09 & ((x10 & ~x11 & x13) | (~x13 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15) | (x07 & (~x11 | (x06 & x11))))))) | (~x10 & ((~x09 & x11 & ((~x06 & (x07 ? (x13 & x16) : (~x13 & ~x16))) | (x07 & x13 & ~x16))) | (~x06 & ~x07 & ~x11 & ~x13))) | (x07 & ~x09 & ~x13))) | (~x13 & ((x08 & ((~x06 & ~x07 & ~x10) | (x09 & x10 & ~x11 & ~x15) | (x07 & (x09 ? ((~x10 & ~x11) | (x06 & (x10 | (~x10 & x11)))) : x11)))) | (~x09 & ((~x06 & ~x07 & x10) | (x07 & ~x11))) | (x09 & x10 & x11 & ~x15))) | (~x11 & x13 & ~x15 & (~x10 | (~x09 & x10)))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x02 & (x04 ? x03 : ~x00)) | (~x00 & x02 & x03 & ~x04 & ((~x08 & ~x09 & ~x10 & x11 & x13) | (~x12 & ~x13 & ((~x09 & ~x10 & x11 & ~x06 & ~x07 & ~x08) | (~x11 & ((x08 & x09 & x10) | (~x06 & ~x07 & ~x08 & (x09 | (~x09 & x10))))))))))))) | (~x00 & x02 & ((x01 & x04) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x04 & ~x06 & ~x07 & ~x01 & x03))) | (~x05 & (x04 ? ((x03 & ((x01 & (x00 ? (x02 & ~x25) : ~x02)) | (x00 & (~x02 | (~x01 & x02))))) | (x00 & ~x01 & ~x03)) : (x02 ? ((~x03 & ((~x12 & ~x13 & ((~x06 & ~x07 & ((((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)) & (x00 | (~x00 & x01))) | (~x08 & x09 & ~x11 & (x01 | (x00 & ~x01))))) | (x08 & x09 & x10 & ~x11 & (x01 | (x00 & ~x01))))) | (~x09 & ~x10 & x11 & x00 & ~x01 & ~x08))) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & x00 & ~x01 & x03 & ~x06 & ~x07)) : (x03 & ~x12 & ~x13 & ((x09 & x10 & ~x11 & ~x01 & x08) | (~x06 & ~x07 & ((x09 & (x08 ? (~x10 & x11) : ~x11) & (~x01 | (~x00 & x01))) | (~x09 & x10 & ~x11 & ~x00 & ~x01 & ~x08)))))))))));
  assign z31 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & ((x05 & ((~x03 & (x00 ? (x01 & (x02 | (~x02 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))))) : ((x02 & ~x04) | (x01 & ~x02 & x04)))) | (x01 & x03 & ((x02 & (~x04 | (x00 & x04))) | (x00 & ~x02 & ~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))))) | (~x01 & ((~x03 & (x00 ? (~x02 | (x02 & x04)) : (x04 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))) | (~x12 & ((~x08 & ((x09 & ((x10 & ~x11 & x13) | (~x13 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15) | (x07 & (~x11 | (x06 & x11))))))) | (~x10 & ((~x09 & x11 & ((~x06 & (x07 ? (x13 & x16) : (~x13 & ~x16))) | (x07 & x13 & ~x16))) | (~x06 & ~x07 & ~x11 & ~x13))) | (x07 & ~x09 & ~x13))) | (~x13 & ((x08 & ((~x06 & ~x07 & ~x10) | (x09 & x10 & ~x11 & ~x15) | (x07 & (x09 ? ((~x10 & ~x11) | (x06 & (x10 | (~x10 & x11)))) : x11)))) | (~x09 & ((~x06 & ~x07 & x10) | (x07 & ~x11))) | (x09 & x10 & x11 & ~x15))) | (~x11 & x13 & ~x15 & (~x10 | (~x09 & x10)))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x02 & (x04 ? x03 : ~x00)) | (~x00 & x02 & x03 & ~x04 & ((~x08 & ~x09 & ~x10 & x11 & x13) | (~x12 & ~x13 & ((~x09 & ~x10 & x11 & ~x06 & ~x07 & ~x08) | (~x11 & ((x08 & x09 & x10) | (~x06 & ~x07 & ~x08 & (x09 | (~x09 & x10))))))))))))) | (~x00 & x02 & ((x01 & x04) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x04 & ~x06 & ~x07 & ~x01 & x03))) | (~x05 & (x04 ? ((x03 & ((x01 & (x00 ? (x02 & ~x25) : ~x02)) | (x00 & (~x02 | (~x01 & x02))))) | (x00 & ~x01 & ~x03)) : (x02 ? ((~x03 & ((~x12 & ~x13 & ((~x06 & ~x07 & ((((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)) & (x00 | (~x00 & x01))) | (~x08 & x09 & ~x11 & (x01 | (x00 & ~x01))))) | (x08 & x09 & x10 & ~x11 & (x01 | (x00 & ~x01))))) | (~x09 & ~x10 & x11 & x00 & ~x01 & ~x08))) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & x00 & ~x01 & x03 & ~x06 & ~x07)) : (x03 & ~x12 & ~x13 & ((x09 & x10 & ~x11 & ~x01 & x08) | (~x06 & ~x07 & ((x09 & (x08 ? (~x10 & x11) : ~x11) & (~x01 | (~x00 & x01))) | (~x09 & x10 & ~x11 & ~x00 & ~x01 & ~x08)))))))))));
  assign z32 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & (x05 ? ((~x03 & (x04 ? (x01 ? (~x02 & x15 & (~x00 | (x00 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (x00 ? (x02 | (~x02 & x15)) : ((x12 & ((~x02 & ~x08 & x09 & ~x10 & ~x11 & x13) | (x02 & ~x06 & ~x07 & ~x13 & x16 & ~x17))) | (x02 & (x17 | (~x17 & ((x13 & (x06 | x15)) | (~x12 & ((~x13 & ((x09 & ((x15 & (x10 | (~x08 & ~x10 & x11))) | (x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10 & x11))))) | (~x06 & ~x07 & ((x08 & ~x10 & x15) | (~x09 & ((x10 & (x08 ? (~x16 & (~x11 | (x11 & x15))) : (~x11 & x15))) | (~x08 & ~x10 & x11 & x15 & ~x16))))))) | (~x08 & ~x09 & ~x06 & x07 & ~x10 & x11 & x13 & x16))))))) | (~x02 & ~x12 & (x13 | (x09 & x11 & ~x13 & (x10 | (~x08 & ~x10)))))))) : (x02 ? (x01 | (~x00 & ~x01)) : x00))) | (~x00 & ~x01 & ~x02 & ~x04) | (x03 & (x02 ? (x01 | (~x00 & ~x01 & ~x04 & ~x06 & ~x07 & ~x11 & ~x12 & ~x13 & ~x08 & x09 & x10)) : ((x00 & ((~x09 & ~x10 & x11 & ~x12 & ~x13 & x15 & ~x06 & ~x07 & ~x08 & x01 & ~x04) | (~x01 & x04 & ~x22))) | (~x00 & ~x01 & x04 & x15))))) : (x01 ? ((x03 & x04 & (~x00 | (x00 & x02 & x25))) | (~x00 & x02 & ~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x08 & x10 & ~x11 & (~x09 | (x09 & x15 & x17))) | (x08 & x09 & ~x10 & x11 & x15)))) : ((~x04 & ((~x00 & ((~x02 & ~x03) | (x11 & ~x12 & ~x13 & x09 & ~x10 & x02 & x03 & ~x06 & ~x07 & x08))) | (~x11 & ~x12 & ~x13 & ~x08 & ~x09 & x10 & x00 & x02 & ~x03 & ~x06 & ~x07))) | (x00 & x04 & (~x02 | (x02 & x03)))))))));
  assign z33 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & ((~x10 & ((~x08 & ((x09 & ((~x02 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (x02 & x11 & ~x12 & ~x13 & ~x17))) | (x02 & ~x09 & ~x17 & ((~x12 & ((x11 & ((~x06 & (x07 ? (x13 & x16) : (~x13 & ~x16))) | (x07 & x13 & ~x16))) | (~x06 & ~x07 & ~x11 & ~x13))) | (x13 & ((x07 & x12) | (x11 & ~x15 & ~x16))))))) | (x02 & ~x17 & ((x08 & ((~x12 & ~x13 & ((~x06 & ~x07 & (x15 | (~x11 & ~x15))) | (x07 & (x09 | (~x09 & x11))))) | (~x09 & x11 & x13 & ~x15))) | (x13 & ~x15 & ((x09 & (x11 | (~x11 & x12))) | (~x11 & ~x12))))))) | (~x12 & (x02 ? (~x17 & ((~x13 & ((x07 & (x09 ? ((x06 & (x08 ? x10 : x11)) | (~x08 & ~x11)) : (~x08 | ~x11))) | (x10 & ((~x06 & ~x07 & ~x09 & (x08 ? (~x16 & (~x11 | (x11 & x15))) : (~x11 & x15))) | (x09 & (x15 | (x11 & ~x15))))))) | (x10 & ~x11 & x13 & (x09 ? ~x08 : ~x15)))) : (x13 | (x09 & x10 & x11 & ~x13)))) | (x02 & (x17 | (~x17 & ((x06 & (~x07 | x13)) | (x13 & ((x10 & (x11 ? ~x15 : ((x12 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (x08 & x09 & ~x15)))) | x15 | (x12 & ~x15 & ~x09 & ~x11))))))))))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((x10 & ~x11 & ~x08 & ~x09) | (x08 & x09 & ~x10 & x11 & x15)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04))))))))));
  assign z34 = x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x00 & ~x01 & x03 & x05) | (~x00 & x01 & ~x02 & (x03 ^ ~x05)))) | (~x20 & ~x21 & (x05 ? ((~x00 & (x04 ? (x01 ? (x02 | (~x02 & ~x03)) : (~x03 & (x02 ? (x17 | (~x17 & ((x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x07 & (x09 ? ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11)) : (~x08 | ~x11 | (x08 & x11)))) | (x10 & ((~x06 & ~x07 & (x08 ? (~x09 & (x16 | (~x16 & (~x11 | (x11 & ~x15))))) : (x11 ? ~x09 : ~x15))) | (x09 & ~x15 & (x11 | (x08 & ~x11))))) | (~x10 & ((~x08 & ((x09 & x11 & ~x15) | (~x06 & ~x07 & (~x11 | (~x09 & x11 & ~x15 & ~x16))))) | (~x06 & ~x07 & x08 & ~x15))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))) : ((x02 & ~x03) | (~x01 & (~x02 | (x02 & x03 & ((~x08 & ~x09 & ~x10 & x11 & x13) | (~x12 & ~x13 & ((x09 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))) | (~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11))))))))))) | (x00 & ((~x03 & (x01 ? (x02 | (~x02 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))))) : (~x02 | (x02 & x04)))) | (x01 & x03 & (x02 ? x04 : (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))))))) | (x03 & (x01 ? (x02 & ~x04) : (~x02 & x04)))) : ((x00 & (x04 ? (~x01 | (x01 & x02 & x03 & ~x25)) : ((~x12 & ~x13 & ((x09 & ((~x01 & ((~x11 & (x02 ^ x03) & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (x02 & x03 & ~x06 & ~x10 & x11 & ~x07 & x08))) | (~x10 & x11 & ~x07 & x08 & x02 & ~x03 & ~x06))) | (x10 & ~x11 & ~x08 & ~x09 & ~x06 & ~x07 & x02 & ~x03))) | (~x10 & x11 & ~x08 & ~x09 & ~x01 & x02 & ~x03)))) | (~x04 & ~x12 & ~x13 & ((~x06 & ~x07 & ((~x02 & x03 & ((~x01 & x08 & x09 & ~x10 & x11) | (~x00 & ((x01 & x09 & (x08 ? (~x10 & x11) : ~x11)) | (~x09 & x10 & ~x11 & ~x01 & ~x08))))) | (x01 & x02 & ~x03 & ((~x08 & x09 & ~x11) | (~x00 & ((x10 & ~x11 & ~x08 & ~x09) | (x08 & x09 & ~x10 & x11 & ~x15))))))) | (x10 & ~x11 & x08 & x09 & x01 & x02 & ~x03))) | (~x00 & x01 & ~x02 & x03 & x04)))));
  assign z35 = ~x14 | (x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((~x01 & ((~x00 & ((~x03 & (x02 ? (x04 & x05 & ((~x17 & ((x07 & (x12 ? ((x13 & ((~x08 & (x09 ? (x10 & ~x11) : ~x10)) | (x10 & ~x11 & x08 & ~x09))) | (x06 & (~x13 | (~x08 & ~x09 & x10 & ~x11 & x13 & ~x15 & x16)))) : ((~x13 & ((x08 & (x09 ? ~x10 : x11)) | (~x09 & ~x11) | (~x08 & (~x09 | (x09 & ~x11))))) | (~x08 & ~x09 & ~x10 & x11 & x13 & (~x16 | (~x06 & x16)))))) | (~x12 & ((~x08 & ((~x13 & ((x09 & ((~x06 & ~x07 & x10 & ~x11 & ~x15) | (~x10 & x11 & x15))) | (~x06 & ~x07 & ((~x10 & ~x11) | (~x09 & (x10 | (~x10 & x11 & ~x16))))))) | (~x11 & x13 & (x09 ? x10 : (~x10 & ~x15))))) | (~x13 & ((~x06 & ~x07 & x08 & ((x15 & (~x10 | (x11 & ~x16 & ~x09 & x10))) | (~x09 & x10 & (x16 | (~x11 & ~x16))))) | (x09 & x10 & x15))))) | (x06 & ~x07) | (~x06 & x12 & ~x13) | (x13 & x15))) | (~x08 & ~x09 & ~x10 & x11 & ~x12 & x16 & x17 & ((x13 & x15) | (~x06 & ~x07 & ~x13 & (~x18 | (x15 & x18))))))) : (x04 ? (x05 & ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))) : (~x05 & (~x25 | (x25 & (~x24 | (x15 & x24)))))))) | (~x02 & ~x04 & x05) | (x03 & (x02 ? (~x04 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : ((~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x06 & ~x07 & ~x08 & ~x04 & ~x05) | (x04 & x05 & x15)))))) | (~x05 & ((x00 & ((~x03 & x04) | (x02 & (x03 ? (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06)) : (~x04 & ((~x11 & ~x12 & ~x13 & x08 & x09 & x10) | (~x08 & ((~x09 & ~x10 & x11) | (~x11 & ~x12 & ~x13 & ~x06 & ~x07 & x09))))))))) | (~x02 & x03 & ~x04 & x09 & ~x12 & ~x13 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))))) | (x00 & x04 & x05 & (x02 ? ~x03 : (x03 | (~x03 & x15)))))) | (x01 & ((~x04 & ((~x12 & ~x13 & (x02 ? (~x03 & ~x05 & ((~x00 & ~x06 & ~x07 & x10 & ~x11 & ~x08 & ~x09) | (x09 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & ((~x00 & x15 & ((x08 & ~x10 & x11) | (~x08 & x10 & ~x11 & x17))) | (~x08 & ~x11 & (~x10 | (x00 & x10))))))))) : (x03 & (x00 ? (x05 & (x09 | (~x06 & ~x07 & ~x08 & ~x09 & ~x10 & x11 & x15))) : (~x05 & ~x06 & ~x07 & x09 & (x08 ? (~x10 & x11) : ~x11)))))) | (x03 & x05 & (x02 | (~x09 & ~x10 & x11 & x13 & x00 & ~x02 & ~x08))))) | (x04 & (x02 ? (~x00 | (x00 & x03)) : (x00 ? (~x03 & x05 & ((x13 & x15) | (x10 & ((~x12 & ~x13 & x15 & x09 & x11) | (~x08 & ~x09 & x06 & x07 & ~x11 & x12 & x13 & ~x15 & x16))))) : (x03 ? ~x05 : (x05 & x15))))) | (x00 & x02 & ~x03 & x05))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ((~x03 & ~x04 & (x02 ? (~x05 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : x05)) | (~x02 & x03 & x04 & ~x05)))))));
  assign z36 = x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x06 & (x13 | (x07 & x12 & ~x13))) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (~x08 & ((x11 & ~x16 & ~x09 & ~x10) | (x09 & x10 & ~x11 & x12))) | (x09 & ~x10) | (x10 & x11) | (~x09 & ~x11 & x12))) | (~x06 & x12 & ~x13) | (~x12 & ((~x09 & x13 & (x10 ? (~x11 & ~x15) : ((x08 & ~x11 & ~x15) | (~x06 & x07 & ~x08 & x11 & x16)))) | (~x13 & ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10 & x11))) | (x10 & ~x15 & (x11 | (x08 & ~x11))) | (~x08 & ~x10 & ((x11 & ~x15) | (~x06 & ~x07 & ~x11))))) | (~x09 & x10 & x11 & x07 & x08) | (~x06 & ~x07 & ((~x15 & (x08 ? (~x10 | (x11 & ~x16 & ~x09 & x10)) : ((x10 & ~x11) | (x11 & ~x16 & ~x09 & ~x10)))) | (~x09 & x10 & (x08 ? (x16 | (~x11 & ~x16)) : x11))))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (x01 & (x02 ? ((~x03 & ((x00 & x05) | (~x04 & ~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))))))))) | (~x00 & x04) | (x03 & ((~x04 & x05) | (x00 & x04 & (x05 | (~x05 & ~x25)))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))))));
  assign z37 = ~x14 | (x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((x02 & ((~x01 & (x00 ? ((~x03 & x04 & x05) | (~x05 & (x03 ? (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06)) : (~x04 & ((~x11 & ~x12 & ~x13 & x08 & x09 & x10) | (~x08 & ((~x09 & ~x10 & x11) | (~x11 & ~x12 & ~x13 & ~x06 & ~x07 & x09)))))))) : ((x11 & ~x12 & ~x13 & x09 & ~x10 & ~x06 & ~x07 & x08 & x03 & ~x04) | (x05 & (x03 ? (~x04 & ((~x08 & ~x09 & ~x10 & x11 & x13) | (~x12 & ~x13 & ((~x09 & ~x10 & x11 & ~x06 & ~x07 & ~x08) | (~x11 & ((x08 & x09 & x10) | (~x06 & ~x07 & ~x08 & (x09 | (~x09 & x10))))))))) : (x04 & (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))))))))) | (x01 & ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))))))))))) | (~x03 & ~x04 & (x00 ? (~x05 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : x05)))) | (x00 & ~x01 & ~x03 & x04 & ~x05) | (~x02 & ((x03 & (x05 ? ((x00 & x01 & ~x04 & ~x12 & ~x13 & (x09 | (~x06 & ~x07 & ~x08 & ~x09 & (x10 ? ~x11 : (x11 & x15))))) | (~x01 & x04)) : (x04 ? (x00 | (~x00 & x01)) : (~x12 & ~x13 & ((~x06 & ~x07 & ((x09 & (x08 ? (~x10 & x11) : ~x11) & (~x01 | (~x00 & x01))) | (~x09 & x10 & ~x11 & ~x00 & ~x01 & ~x08))) | (x09 & x10 & ~x11 & ~x00 & ~x01 & x08)))))) | (~x01 & (x00 ? (~x03 & x05) : (~x04 & (x05 | (~x03 & ~x05))))) | (x00 & x01 & ~x03 & x05 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))))))))));
  assign z38 = ~x14 | (x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (x08 & ~x09 & ~x10 & ~x11 & ~x15)) : ((x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11) | (x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (x10 & (x15 | (x08 & ~x11 & ~x15))) | (~x08 & ((~x06 & ~x07 & x10 & ~x11 & ~x15) | (~x10 & x11 & x15)))))))) | (x13 & ((x12 & ((~x09 & ~x10 & x07 & ~x08) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x15 & (~x09 | (x08 & x09 & ~x10))))))) | x06 | x15 | (~x08 & ~x09 & ~x10 & x11 & ~x15 & ~x16))) | (~x06 & x12 & ~x13) | (x06 & (~x07 | (x07 & x12 & ~x13)))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z39 = ~x14 | (x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((x05 & (x02 ? (x03 ? ((x01 & ~x04) | (~x00 & ((~x13 & ((~x06 & ~x07 & (x01 ? (x04 & x16 & (x12 | (x08 & ~x09 & x10 & x11 & ~x12))) : (~x04 & ~x08 & ~x12 & (x09 ? ~x11 : (x10 ^ x11))))) | (~x01 & ~x04 & x08 & x09 & x10 & ~x11 & ~x12))) | (~x09 & ~x10 & x11 & x13 & ~x01 & ~x04 & ~x08)))) : ((x00 & (x01 ? (~x04 & ~x24) : x04)) | (x01 & x04) | (~x00 & ~x01 & (x04 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (x12 & (x13 ? ((~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15))) | (~x09 & ~x10 & x07 & ~x08)) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x10 & x11) | (~x10 & (x09 | (x11 & ~x16 & ~x08 & ~x09))))) | (~x12 & (x13 ? ((~x09 & (x10 ? (~x11 & ~x15) : ((x08 & ~x11 & ~x15) | (x07 & ~x08 & x11 & (~x16 | (~x06 & x16)))))) | (x10 & ~x11 & ~x08 & x09)) : ((x09 & ((~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))) | (x07 & ((x06 & (x08 ? x10 : x11)) | (~x08 & ~x11) | (x08 & ~x10 & (~x11 | (~x06 & x11))))))) | (~x09 & (((x07 | (~x06 & ~x07 & x10)) & (~x08 | (x08 & x11))) | (x07 & ~x11) | (~x06 & ~x07 & ~x08 & ~x10 & x11 & ~x16))) | (~x06 & ~x07 & ~x10 & (x08 | (~x08 & ~x11))))))))) : ~x23)))) : (x00 ? (x01 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 | (x03 & x04 & x22))) : ((~x01 & x03) | (x04 & x15 & x01 & ~x03))))) | (x03 & ~x04 & ~x06 & ~x00 & ~x01 & x02 & ~x07 & x08 & x09 & ~x12 & ~x13 & ~x10 & x11) | (~x05 & (x04 ? ((~x00 & x01 & ~x02 & x03) | (x00 & (~x01 | (x01 & x02 & x03)))) : ((~x12 & ~x13 & ((~x06 & ~x07 & (x02 ? (~x03 & ((((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)) & (x00 | (~x00 & x01))) | (~x08 & x09 & ~x11 & (x01 | (x00 & ~x01))))) : (x03 & x09 & ((~x10 & ((~x01 & (x08 ^ ~x11)) | (x08 & x11 & ~x00 & x01))) | (~x08 & x10 & ~x11 & x00 & ~x01))))) | (x08 & x09 & x10 & ~x11 & (x01 ? (x02 & ~x03) : (x00 ? (x02 & ~x03) : (~x02 & x03)))))) | (~x00 & ~x01 & ~x02 & ~x03 & (~x25 | (~x15 & x24 & x25))))))))));
  assign z40 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (((~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)) & (x02 ^ ~x05)) | (~x02 & x05) | (x02 & x03 & ((x05 & ~x08 & ~x09 & ~x10 & x11 & x13) | (~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (~x10 & x11 & ~x08 & ~x09 & x05 & ~x06 & ~x07))))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (~x06 & ~x07 & ~x10 & (x08 | (~x08 & ~x11))) | (~x09 & ((x11 & ((~x06 & ~x07 & ~x16 & (~x08 ^ x10)) | (x07 & x08 & ~x10))) | (x07 & (~x08 | ~x11)) | (~x06 & ~x07 & x10 & ~x11)))))) | (x06 & (~x07 | x13)) | (~x06 & ~x07 & x12 & ~x13) | (x13 & ((~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))) | (x12 & ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))))) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (x01 & (x02 ? (x04 ? (~x00 | (x00 & (x03 ? (x05 | (~x05 & x25)) : (x05 & ~x16)))) : (x05 | (~x03 & ~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04))))))))));
  assign z41 = ~x14 | (x14 & ((~x19 & (x20 | x21)) | (~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x20 & ~x21 & ((x05 & ((~x00 & (x04 ? (x01 ? (x02 | (~x02 & ~x03)) : (~x03 & (x02 ? (x17 | (~x17 & ((~x12 & (x13 ? ((~x09 & (x10 ? (~x11 & ~x15) : ((x08 & ~x11 & ~x15) | (x07 & ~x08 & x11 & (~x16 | (~x06 & x16)))))) | (x10 & ~x11 & ~x08 & x09)) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & (x15 | (~x15 & (x11 | (x08 & ~x11))))))) | (x08 & ~x10 & ~x06 & ~x07) | (~x09 & ((x08 & ((~x06 & ~x07 & x10) | (x07 & x11))) | (x07 & (~x08 | ~x11)) | (~x06 & ~x07 & ~x08 & (x10 ? (x11 | (~x11 & x15)) : (~x11 | (x11 & ~x16))))))))) | (x12 & (x13 ? ((~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15))) | (~x09 & ~x10 & x07 & ~x08)) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & (x15 | (~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x10 & x11) | (~x10 & (x09 | (x11 & ~x16 & ~x08 & ~x09)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))) : ((x02 & ~x03) | (~x01 & (~x02 | (x02 & x03 & ~x12 & ~x13 & ((~x09 & ~x10 & x11 & ~x06 & ~x07 & ~x08) | (~x11 & ((x08 & x09 & x10) | (~x06 & ~x07 & ~x08 & (x09 | (~x09 & x10)))))))))))) | (x03 & (x01 ? (x02 & ~x04) : (~x02 & x04))) | (x00 & ((~x03 & (x01 ? (x02 | (~x02 & (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13)))))) : (~x02 | (x02 & x04)))) | (x01 & ~x02 & x03 & ~x04 & ~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))))) | (~x05 & (x04 ? (x00 ? ~x01 : (x01 & x03)) : (x00 ? (x02 & ~x03 & ~x12 & ~x13 & ((~x01 & ~x06 & ~x07 & ((~x08 & x10 & ~x11) | (~x10 & x11 & x08 & x09))) | (x09 & x10 & ~x11 & x01 & x08))) : (x01 ? (~x06 & ~x07 & ~x12 & ~x13 & ((~x09 & x10 & ~x11 & x02 & ~x03 & ~x08) | (x09 & ((~x02 & x03 & x08 & ~x10 & x11) | (x02 & ~x03 & (x08 ? (~x10 & x11) : ~x11)))))) : ((~x02 & ~x03) | (x11 & ~x12 & ~x13 & x09 & ~x10 & x02 & x03 & ~x06 & ~x07 & x08)))))) | (x00 & x01 & x02 & x03 & x04)))));
  assign z42 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & (x05 ? ((~x03 & (x00 ? (~x02 | (x02 & x04)) : (x04 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (~x02 & (x04 ? x03 : ~x00)) | (~x00 & x02 & x03 & ~x04 & ((~x12 & ~x13 & ((x09 & ((~x06 & ~x07 & ~x10 & (x08 ^ ~x11)) | (x08 & x10 & ~x11))) | (~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (~x08 & ~x09 & ~x10 & x11 & x13)))) : ((~x04 & ((~x02 & ((~x00 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06))) | (x03 & x09 & ~x12 & ~x13 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))))) | (x00 & x02 & ((x09 & ~x12 & ~x13 & ((~x03 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (x08 & ~x10 & x11 & x03 & ~x06 & ~x07))) | (~x09 & ~x10 & x11 & ~x03 & ~x08))))) | (x00 & x04 & (~x03 | (x02 & x03)))))) | (x01 & ((x00 & ((~x04 & ((~x08 & ((~x06 & ~x07 & ~x12 & ~x13 & ((~x11 & ((x02 & ~x03 & ~x05 & (x10 | (x09 & ~x10))) | (~x02 & x03 & x05 & ~x09 & x10))) | (~x09 & ~x10 & x11 & ~x02 & x03 & x05))) | (~x09 & ~x10 & x11 & x13 & ~x02 & x03 & x05))) | (~x02 & x05 & (~x03 | (~x12 & ~x13 & x03 & x09))))) | (x02 & (x03 ? x04 : x05)) | (~x02 & ~x03 & x04 & x05 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) | (x05 & ((~x00 & ~x02 & ~x03 & x04) | (x02 & x03 & ~x04))) | (~x00 & (x04 ? (x02 | (~x02 & x03 & ~x05)) : (~x05 & ~x06 & ~x07 & ~x12 & ~x13 & ((x09 & (x02 ^ x03) & (x08 ? (~x10 & x11) : ~x11)) | (~x09 & x10 & ~x11 & x02 & ~x03 & ~x08))))) | (x09 & x10 & ~x11 & ~x12 & ~x13 & x02 & ~x03 & ~x04 & ~x05 & x08))) | (x00 & ~x05 & ((~x02 & x03 & x04) | (x02 & ~x03 & ~x04 & ~x06 & ~x07 & x11 & ~x12 & ~x13 & x08 & x09 & ~x10))) | (~x00 & x02 & ~x03 & ~x04 & x05)))));
  assign z43 = x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & ((~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))) | (((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & ~x02 & x03 & ~x04) | (x00 & ((~x05 & ((~x03 & x04) | (x02 & ~x04 & ~x10 & x11 & ((~x03 & ~x08 & ~x09) | (x03 & ~x06 & ~x07 & ~x12 & ~x13 & x08 & x09))))) | (~x02 & ~x03 & x05))))) | (x01 & (x02 ? ((x05 & (x03 ? ~x04 : x00)) | (~x00 & x04) | (~x03 & ~x04 & ~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & ((x03 & x04) | (x02 & ~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))))))));
  assign z44 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z45 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z46 = x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))) | (~x04 & ((~x02 & ~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06))) | (~x03 & x05) | (x02 & x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))))))))) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (x01 & (x02 ? ((x00 & (x03 ? (x04 & (x05 | (~x05 & ~x25))) : x05)) | (~x00 & x05) | (~x05 & ((~x00 & x04) | (~x03 & ~x04 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))))));
  assign z47 = x14 & ((~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((~x00 & ((~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))) | (~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06))))))) | (~x02 & ((x05 & (x03 ^ ~x04)) | (x03 & ~x04 & ~x05 & x09 & ~x12 & ~x13 & ((x08 & x10 & ~x11) | (~x06 & ~x07 & (x08 ? (~x10 & x11) : ~x11)))))) | (x00 & ((~x03 & x04) | (x02 & ~x05 & (x03 ? (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06)) : (~x04 & ((~x11 & ~x12 & ~x13 & x08 & x09 & x10) | (~x08 & ((~x09 & ~x10 & x11) | (~x11 & ~x12 & ~x13 & ~x06 & ~x07 & x09))))))))))))) | (~x19 & (x20 | x21)) | (~x04 & x05 & (x00 ? (~x01 & (x02 ^ x03)) : (x01 & ~x02))));
  assign z48 = ~x14 | (x14 & ((~x03 & ~x04 & x05 & (x00 ? (~x01 & x02) : (x01 & ~x02))) | (~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z49 = ~x14 | (x14 & ((~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))))))) | (~x04 & ((~x00 & x01 & ~x02 & ~x03) | (x00 & ~x01 & x05 & (x02 ^ x03)))) | (~x19 & (x20 | x21))));
  assign z50 = ~x14 | (x14 & ((~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))))))))) | (~x04 & ((~x00 & x01 & ~x02 & ~x03) | (x00 & ~x01 & x05 & (x02 ^ x03)))) | (~x19 & (x20 | x21))));
  assign z51 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((x01 & (x02 ? ((x00 & (x03 ? x04 : x05)) | (~x00 & x04) | (~x04 & (x03 ? x05 : (~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & (x02 ? (~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))) : (x03 & x04))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (~x02 & ((x00 & ~x03 & x05) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & x03 & ~x04))) | (x00 & ~x05 & ((~x03 & x04) | (x02 & ((x03 & (x04 | (x11 & ~x12 & ~x13 & x09 & ~x10 & ~x07 & x08 & ~x04 & ~x06))) | (~x09 & ~x10 & x11 & ~x03 & ~x04 & ~x08))))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x05 | (~x05 & (~x03 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & x03 & ~x06)))))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (~x11 & ((x07 & ~x09) | (~x06 & ~x07 & ~x08 & ~x10))) | (x08 & ~x10 & ~x06 & ~x07) | (~x09 & ((x07 & (~x08 | (x08 & x11))) | (~x06 & ~x07 & ((~x08 & ~x10 & x11 & ~x16) | (x10 & (~x08 | (x08 & (x16 | (x11 & ~x16))))))))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z52 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((x01 & (x02 ? ((x05 & (x03 ? ~x04 : x00)) | (~x00 & x04) | (~x03 & ~x04 & ~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (~x00 & x02 & ~x03 & ~x04 & x05) | (x00 & ~x05 & ((x03 & x04) | (x02 & ~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09))))) | (~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & ~x02 & x03 & ~x04) | (x00 & ((~x05 & ((~x03 & x04) | (x02 & ~x04 & ~x10 & x11 & ((~x03 & ~x08 & ~x09) | (x03 & ~x06 & ~x07 & ~x12 & ~x13 & x08 & x09))))) | (~x02 & ~x03 & x05))) | (~x00 & ((~x04 & (x02 ? (x03 & ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13))) : (x03 ? (x05 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & ~x05 & ~x06)) : ~x05))) | (~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16))))))) | (~x12 & ((~x08 & ((x09 & ((x10 & ~x11 & x13) | (~x13 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15) | (x07 & (~x11 | (x06 & x11))))))) | (~x10 & ((~x09 & x11 & ((~x06 & (x07 ? (x13 & x16) : (~x13 & ~x16))) | (x07 & x13 & ~x16))) | (~x06 & ~x07 & ~x11 & ~x13))) | (x07 & ~x09 & ~x13))) | (~x11 & x13 & ~x15 & (~x10 | (~x09 & x10))) | (~x13 & ((~x09 & ((~x06 & ~x07 & x10) | (x07 & ~x11))) | (x09 & x10 & x11 & ~x15) | (x08 & ((~x06 & ~x07 & ~x10) | (x09 & x10 & ~x11 & ~x15) | (x07 & (x09 ? ((~x10 & (~x11 | (~x06 & x11))) | (x06 & (x10 | (~x10 & x11 & x18)))) : x11))))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11))))))))))))));
  assign z53 = ~x14 | (x14 & ((~x04 & ((x05 & ((x00 & ~x01 & (x02 | (~x02 & x03))) | (~x00 & x01 & ~x02 & x03))) | (~x00 & x01 & ~x02 & ~x03))) | (~x19 & (x20 | x21)) | (~x20 & ~x21 & ((~x01 & ((((~x02 & x03) | (x00 & x02 & ~x03)) & (x04 ? x05 : (~x05 & x09 & ~x11 & ~x12 & ~x13 & ((x08 & x10) | (~x06 & ~x07 & ~x08))))) | (x11 & ~x12 & ~x13 & x08 & x09 & ~x10 & ~x05 & ~x06 & ~x07 & ~x02 & x03 & ~x04) | (x00 & ((~x05 & ((~x03 & x04) | (x02 & ~x04 & ~x10 & x11 & ((~x03 & ~x08 & ~x09) | (x03 & ~x06 & ~x07 & ~x12 & ~x13 & x08 & x09))))) | (~x02 & ~x03 & x05))) | (~x00 & ((~x03 & x04 & x05 & (x02 ? (x17 | (~x17 & ((x15 & (x13 | (x09 & x10 & ~x12 & ~x13))) | (~x12 & (x13 ? ((~x08 & ((x07 & ~x09 & ~x10 & x11 & (~x16 | (~x06 & x16))) | (x09 & x10 & ~x11))) | (~x11 & ~x15 & (~x10 | (~x09 & x10)))) : ((x09 & ((x07 & ((x06 & (x08 ? x10 : x11)) | (x08 & ~x10) | (~x08 & ~x11))) | (~x08 & ((~x10 & x11) | (~x06 & ~x07 & x10 & ~x11 & ~x15))) | (x10 & ~x15 & (x11 | (x08 & ~x11))))) | (x08 & ((~x06 & ~x07 & ~x10) | (x07 & ~x09 & x11))) | (~x09 & ((~x06 & ~x07 & (x10 | (~x08 & ~x10 & x11 & ~x16))) | (x07 & (~x08 | ~x11)))) | (~x06 & ~x07 & ~x08 & ~x10 & ~x11)))) | (x12 & (x13 ? ((~x10 & ((x07 & ~x08 & ~x09) | (x09 & ~x11 & ~x15))) | (~x11 & ((x10 & ((x07 & (x08 ^ x09)) | (~x08 & x09 & ~x15))) | (~x09 & ~x15)))) : (~x06 | (x06 & x07)))) | (x06 & (~x07 | x13)) | (x13 & ~x15 & ((x08 & (x09 ? (x10 & ~x11) : (~x10 & x11))) | (x11 & (x10 | (~x10 & (x09 | (~x08 & ~x09 & ~x16)))))))))) : ((~x12 & x13) | (x09 & ((~x08 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13))) | (~x12 & ~x13 & x10 & x11)))))) | (~x04 & (x03 ? (x02 ? ((~x12 & ~x13 & ((x09 & ((x05 & ~x11 & ((x08 & x10) | (~x06 & ~x07 & ~x08))) | (~x06 & ~x07 & x08 & ~x10 & x11))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & (x10 ^ x11)))) | (x05 & ~x08 & ~x09 & ~x10 & x11 & x13)) : (x05 | (~x09 & x10 & ~x11 & ~x12 & ~x13 & ~x07 & ~x08 & ~x05 & ~x06))) : (x02 ? (x05 & x23) : ~x05))))))) | (x01 & (x02 ? ((x05 & (x03 ? ~x04 : x00)) | (~x00 & x04) | (~x03 & ~x04 & ~x05 & ~x12 & ~x13 & ((x10 & ~x11 & x08 & x09) | (~x06 & ~x07 & ((~x08 & x09 & ~x11) | (~x00 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))) : ((~x00 & x03 & ~x05 & (x04 | (~x04 & ~x06 & ~x07 & x09 & ~x12 & ~x13 & (x08 ? (~x10 & x11) : ~x11)))) | (x05 & (x00 ? (x03 ? (~x04 & ((x09 & ~x12 & ~x13) | (~x08 & ~x09 & ((~x10 & x11 & x13) | (~x06 & ~x07 & ~x12 & ~x13 & (x10 ^ x11)))))) : (~x04 | (x04 & (x13 | (x09 & x10 & x11 & ~x12 & ~x13))))) : (~x03 & x04)))))) | (x00 & ~x05 & ((x03 & x04) | (x02 & ~x03 & ~x04 & ~x06 & ~x07 & ~x12 & ~x13 & ((~x10 & x11 & x08 & x09) | (x10 & ~x11 & ~x08 & ~x09)))))))));
endmodule