module pla__table5 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14;
  assign z00 = x03 & ~x04 & ~x07 & x08 & ~x10 & ~x13 & (x00 ? (x01 & ~x02 & x09 & (x14 | x15)) : (~x01 & x02 & ~x09 & ~x11 & x12 & (x14 | (x15 & x16))));
  assign z01 = (~x13 & (x01 ? ((~x14 & ~x15 & (x00 ? (x06 & ((~x02 & ~x04 & ~x07 & ~x08 & ~x09 & ~x10 & ~x11 & ~x12 & x16) | (x02 & ~x03 & x04 & x05 & x07 & ~x16))) : (~x03 & ~x05 & ~x06 & ~x16 & ((x02 & x04 & x07) | (~x02 & ~x04 & ~x07 & ~x08 & ~x11 & ~x12 & ~x09 & ~x10))))) | (~x00 & x02 & ~x03 & ~x04 & (x14 | x15 | (~x08 & ~x09 & ~x06 & ~x07 & ~x12 & x16 & ~x10 & ~x11)))) : ((~x02 & ((~x07 & ((~x10 & ((x09 & (((x14 | x15) & ((x00 & ~x04 & (~x08 | (x03 & x08 & ~x11 & ~x12))) | (~x00 & x03 & x04 & ~x08))) | (x03 & x04 & ~x08 & ~x14 & x15 & ~x16))) | (x00 & ~x04 & ~x09 & ~x11 & ((~x03 & x08 & (x14 | (x15 & x16))) | (x03 & x06 & ~x08 & ~x12 & ~x14 & ~x15 & x16))))) | (~x00 & x03 & x04 & ((x08 & (x14 | x15)) | (~x08 & x09 & x10 & ~x11 & x15 & ~x16 & x12 & ~x14))))) | (~x00 & x03 & x04 & ~x14 & ~x15 & (x05 ? (x06 & x07 & (x08 | (~x08 & ~x16))) : (~x06 & ~x16))))) | (x00 & ~x07 & ((~x10 & ((~x12 & ((x02 & ((x09 & ((x08 & (x14 | x15) & (x03 ? (x04 & x11) : (~x04 & ~x11))) | (~x03 & x04 & ~x08 & x15 & ~x16 & x11 & ~x14))) | (~x04 & x06 & ~x08 & ~x09 & ~x15 & x16 & ~x11 & ~x14))) | (x06 & ~x08 & ~x03 & ~x04 & ~x09 & ~x11 & ~x14 & ~x15 & x16))) | (x04 & ~x08 & x02 & x03 & ~x14 & x15 & ~x16 & x09 & ~x11))) | (x02 & ~x03 & x04 & ~x08 & ~x09 & ~x14 & x15 & ~x16 & x10 & x11 & x12))) | (~x14 & ~x15 & x16 & ~x00 & x03 & x04)))) | (~x04 & ((x02 & (x00 ? ((x01 & x03) | (~x01 & ~x03 & x05 & x06 & x07 & x13)) : (x01 & x03 & ~x05 & x07 & x13 & (x14 ^ x15)))) | (~x00 & ~x01 & ~x02 & ~x03))) | (~x00 & ~x02 & x04 & ~x05 & x07 & x08 & ~x09 & ~x10 & x13 & ((x14 & ~x15 & (x11 ^ x12) & (x01 ? (~x03 & ~x16) : x03)) | (~x01 & x03 & ~x14 & x15 & x16 & (~x12 | (~x11 & x12)))));
  assign z02 = x02 ? (x03 ? ((~x01 & ((~x04 & ((x00 & ((x07 & x13 & x05 & x06) | (~x07 & ~x08 & x09 & ~x10 & x15 & ~x16 & ~x13 & ~x14))) | (~x00 & x05 & x06 & x07 & ~x13 & ~x14 & ~x15 & ~x16))) | (~x00 & x04 & ~x07 & ~x08 & x09 & x10 & ~x11 & ~x12 & ~x13 & (x14 | x15)))) | (~x00 & x01 & ((x04 & ((~x05 & x07 & ((x13 & (x14 ^ x15)) | (~x06 & ~x13 & ~x14 & ~x15 & ~x16))) | (~x06 & ~x13 & (x14 | x15)))) | (~x04 & ~x06 & ~x07 & ~x08 & ~x09 & ~x10 & ~x14 & ~x15 & x16 & ~x11 & ~x12 & ~x13)))) : (~x13 & ((x04 & (((x14 | x15) & ((~x00 & x01) | (x00 & ~x01 & ~x07 & x08 & ~x11 & ~x12 & x09 & ~x10))) | (~x00 & ~x06 & ~x14 & ~x15 & ((~x12 & x16 & ~x10 & ~x11 & ~x08 & ~x09 & x01 & ~x07) | (~x01 & ~x05 & ~x16))))) | (~x14 & ~x15 & x16 & ~x00 & ~x01 & ~x04)))) : ((~x13 & ((~x07 & ~x11 & ((x03 & ~x12 & ((x09 & (x14 | x15) & ((~x00 & x01 & ~x04 & ~x08 & x10) | (x00 & ~x01 & x04 & x08 & ~x10))) | (~x00 & x01 & ~x04 & ~x05 & ~x06 & ~x14 & ~x15 & ~x16 & ~x08 & ~x09 & ~x10))) | (x00 & x01 & ~x03 & ~x04 & ~x08 & ~x14 & x15 & ~x16 & x09 & ~x10))) | (~x00 & x01 & ~x03 & ~x15 & x16 & ~x04 & ~x14))) | (~x00 & x01 & x03 & x04 & ~x05 & x07 & x08 & x13 & x14 & ~x15));
  assign z03 = (x02 & ((~x03 & (x04 ? (x00 ? ((x07 & ((x05 & x06 & ((~x01 & x13) | (~x14 & ~x15 & ~x16 & x01 & ~x13))) | (x01 & ~x05 & x13 & ((~x09 & ((~x10 & ((x11 & ((x15 & ~x16 & x12 & ~x14) | (x08 & ~x12 & x14 & ~x15 & x16))) | (x08 & ~x11 & x16 & (x12 ? (x14 & ~x15) : (~x14 & x15))))) | (~x14 & x15 & ~x16 & x10 & ~x11 & ~x12))) | (x15 & ~x16 & ~x08 & ~x14))))) | (~x01 & ~x07 & ~x08 & x11 & ~x13 & ~x14 & x15 & ~x16 & (x09 ? (~x10 & ~x12) : (x10 & x12)))) : (~x13 & ((~x14 & ~x15 & ((~x09 & ~x10 & ~x11 & ~x12 & x16 & ~x07 & ~x08 & x01 & ~x06) | (~x01 & x05 & x06 & x07 & ~x16))) | (x01 & (x14 | x15))))) : ((~x13 & (((x14 | x15) & (~x00 | (x00 & ~x01 & ~x07 & x08 & ~x11 & ~x12 & x09 & ~x10))) | (~x00 & ((~x06 & ((~x12 & x16 & ~x10 & ~x11 & ~x08 & ~x09 & x01 & ~x07) | (~x01 & ~x05 & ~x16))) | (~x01 & ((~x14 & ~x15 & x16) | (x07 & ~x16 & x05 & x06))))))) | (~x00 & ~x01 & ~x05 & x07 & x08 & (x14 ? ~x15 : (x15 & x16)))))) | (~x04 & ((~x01 & ((x05 & x06 & x07 & ((x00 & x13) | (~x14 & ~x15 & ~x16 & ~x00 & x03 & ~x13))) | (x03 & ~x13 & ((~x07 & x09 & (((x14 | x15) & ((x00 & x08 & ~x10) | (x10 & ~x11 & ~x12 & ~x00 & ~x08))) | (~x14 & x15 & ~x16 & x00 & ~x08 & ~x10))) | (~x14 & ~x15 & ~x16 & ~x00 & ~x05 & ~x06))))) | (~x00 & x01 & x03 & ((~x14 & ((~x05 & x07 & ((x13 & x15) | (~x15 & ~x16 & ~x06 & ~x13))) | (~x06 & ~x07 & ~x08 & ~x09 & ~x10 & ~x11 & ~x12 & ~x13 & ~x15 & x16))) | (x13 & x14 & ~x15 & ~x05 & x07))))) | (x04 & ((~x14 & ((~x00 & x01 & ~x05 & x07 & ((x13 & x15) | (~x15 & ~x16 & ~x06 & ~x13))) | (~x01 & x03 & ~x07 & ~x08 & ~x10 & ~x11 & ~x13 & ((x06 & ~x09 & ~x12 & ~x15 & x16) | (x15 & ~x16 & x00 & x09))))) | (~x00 & x01 & ~x05 & x07 & x13 & x14 & ~x15))))) | (~x02 & (x01 ? ((~x13 & ((~x14 & ((~x03 & ((~x00 & ~x15 & x16) | (~x07 & ~x08 & x00 & ~x04 & x09 & ~x10 & ~x11 & x15 & ~x16))) | (~x00 & x04 & ~x06 & ~x07 & ~x08 & ~x09 & ~x10 & ~x11 & ~x12 & ~x15 & (x16 ? x03 : ~x05)))) | (~x00 & x03 & ~x07 & ~x08 & x09 & x10 & ~x11 & ~x12 & (x14 | x15)))) | (~x00 & x03 & ~x04 & ~x05 & x07 & x08 & x13 & x14 & ~x15 & ~x16)) : (x00 ? (~x07 & ~x10 & ~x11 & ~x12 & ~x13 & ((x03 & x08 & x09 & (x14 | x15)) | (x06 & ~x08 & ~x03 & x04 & ~x15 & x16 & ~x09 & ~x14))) : (~x03 & x04)))) | (~x13 & ((~x03 & ~x07 & x09 & ~x11 & ~x12 & (x14 | x15) & ((~x00 & x01 & ~x04 & ~x08 & x10) | (x00 & ~x01 & x04 & x08 & ~x10))) | (~x14 & ~x15 & x16 & ~x00 & ~x01 & x03)));
  assign z04 = x02 ? ((x04 & (x01 ? ((~x14 & ((x07 & ((~x05 & (x00 ? (~x03 & x13 & x15 & ((~x08 & ~x16) | (~x09 & ((~x10 & ((~x12 & x16 & x08 & ~x11) | (x11 & x12 & ~x16))) | (x10 & ~x11 & ~x12 & ~x16))))) : (x03 & ((x13 & x15) | (~x15 & ~x16 & ~x06 & ~x13))))) | (x00 & ~x03 & x05 & ~x15 & ~x16 & x06 & ~x13))) | (~x00 & ~x03 & ~x06 & ~x07 & ~x08 & ~x09 & ~x13 & ~x15 & x16 & ~x10 & ~x11 & ~x12))) | (~x05 & x07 & x13 & x14 & ~x15 & (x00 ? (~x03 & x08 & ~x09 & ~x10 & x16 & (x11 ^ x12)) : x03))) : (~x13 & ((~x07 & x09 & ~x11 & ~x12 & (x14 | x15) & ((~x00 & x03 & ~x08 & x10) | (x08 & ~x10 & x00 & ~x03))) | (~x00 & ~x03 & ~x05 & ~x15 & ~x16 & ~x06 & ~x14))))) | (~x01 & ((x03 & (x00 ? ((x07 & x13 & x05 & x06) | (~x08 & x09 & ~x04 & ~x07 & ~x14 & x15 & ~x16 & ~x10 & ~x13)) : (~x04 & ~x13 & ~x14 & ~x15 & ~x16 & (x05 ? (x06 & x07) : ~x06)))) | (~x14 & ~x15 & x16 & ~x00 & ~x03 & ~x13)))) : ((~x13 & ((~x07 & ~x11 & ((x00 & x01 & ~x03 & ~x04 & ~x08 & ~x14 & x15 & ~x16 & x09 & ~x10) | (x03 & ~x12 & ((x09 & (x14 | x15) & ((x00 & ~x01 & x04 & x08 & ~x10) | (~x00 & x01 & ~x08 & x10))) | (~x00 & x01 & ~x05 & ~x06 & ~x08 & ~x09 & ~x10 & ~x14 & ~x15 & ~x16))))) | (~x03 & ~x14 & ~x15 & ((~x00 & x01 & x16) | (x00 & ~x01 & ~x04 & x07 & ~x16 & ~x05 & ~x06))))) | (~x03 & x04 & ~x00 & ~x01));
  assign z05 = (~x13 & ((~x01 & ((~x07 & ((x00 & ((~x03 & ((~x10 & ((~x11 & ((x08 & ((x09 & ~x12 & (x14 | x15) & (x02 ^ x04)) | (~x02 & ~x04 & ~x09 & (x14 | (x15 & x16))))) | (x06 & ~x08 & ~x09 & ~x12 & ~x14 & ~x15 & x16 & (~x04 | (~x02 & x04))))) | (~x08 & x09 & x02 & x04 & ~x14 & x15 & ~x16 & x11 & ~x12))) | (x02 & x04 & ~x08 & ~x09 & x10 & ~x14 & x15 & ~x16 & x11 & x12))) | (~x10 & ((x04 & ~x08 & x02 & x03 & ~x14 & x15 & ~x16 & x09 & ~x11) | (~x04 & ((~x08 & ((~x02 & x09 & (x14 | x15)) | (x06 & ~x09 & ~x11 & ~x12 & ~x14 & ~x15 & x16 & (x02 | (~x02 & x03))))) | (x03 & x08 & x09 & (x14 | x15) & (x02 | (~x02 & ~x11 & ~x12))))))))) | (~x00 & (((x14 | x15) & ((~x08 & x09 & ((x02 & ((~x03 & x04 & ~x10) | (x10 & ~x11 & ~x12 & x03 & ~x04))) | (~x02 & x03 & x04 & ~x10))) | (~x02 & x03 & x04 & x08))) | (x04 & ~x11 & ((x02 & ~x03 & x08 & ~x09 & ~x10 & ~x12 & (x14 | x16)) | (~x08 & x09 & ~x02 & x03 & ~x14 & x15 & ~x16 & x10 & x12))))) | (x03 & x04 & ~x08 & ~x10 & ~x14 & ((x02 & x06 & ~x09 & ~x11 & ~x12 & ~x15 & x16) | (x15 & ~x16 & ~x02 & x09))))) | (~x00 & ((~x16 & ((~x14 & ~x15 & ((x05 & x06 & x07 & ((x02 & (x03 ^ x04)) | (x04 & ~x08 & ~x02 & x03))) | (~x02 & x03 & x04 & ~x05 & ~x06))) | (x02 & ~x03 & ~x04 & (x05 ? (x06 & x07) : ~x06)))) | (~x14 & ~x15 & ((x03 & (x16 | (~x02 & x04 & x05 & x06 & x07 & x08))) | (x02 & ~x03 & x04 & x16))))) | (x00 & ~x02 & ~x03 & ~x04 & ~x05 & ~x14 & ~x15 & ~x16 & ~x06 & x07))) | (~x00 & ((x01 & ((~x06 & (x02 ? (x03 ? ((x04 & (x14 | x15)) | (~x14 & ~x15 & ~x16 & ~x04 & ~x05 & x07)) : ((~x12 & x16 & ~x10 & ~x11 & ~x08 & ~x09 & ~x04 & ~x07) | (~x14 & ~x15 & ~x16 & x04 & ~x05 & x07))) : (~x07 & ~x08 & ~x09 & ~x10 & ~x11 & ~x12 & ~x14 & ~x15 & (x04 ? (x03 ? x16 : (~x05 & ~x16)) : (~x05 & ~x16))))) | (~x03 & ~x04 & ~x07 & ~x08 & x09 & x10 & ~x11 & ~x12 & (x14 | x15)))) | (x02 & ~x03 & ~x04 & (x14 | x15)))) | (x00 & x01 & ~x02 & ~x04 & x06 & ~x07 & ~x08 & ~x12 & ~x14 & ~x15 & x16 & ~x09 & ~x10 & ~x11))) | (x07 & ((x13 & ((~x01 & ((x02 & (x00 ? (x05 & x06 & (x04 | (~x03 & ~x04))) : (x03 & x04 & ~x05 & x08 & (x14 ? ~x15 : (x15 & x16))))) | (~x00 & ~x02 & x03 & x04 & ~x05 & x08 & ~x09 & ~x10 & ((~x11 & x12 & (x14 ? ~x15 : (x15 & x16))) | (~x12 & ((~x14 & x15 & x16) | (x11 & x14 & ~x15))))))) | (~x00 & x01 & ~x05 & (x02 ? ((x14 ^ x15) & (x03 ^ x04)) : ((x08 & ((x14 & ~x15 & (x03 ? (x04 | (~x04 & ~x16)) : (~x04 | (x04 & ~x09 & ~x10 & ~x16 & (x11 ^ x12))))) | (~x03 & ~x04 & ~x14 & x15 & x16))) | (~x14 & x15 & ~x16 & ~x03 & ~x04)))))) | (~x00 & ~x01 & x02 & ~x03 & ~x04 & ~x05 & x08 & (x14 ? ~x15 : (x15 & x16))))) | (~x04 & ((~x00 & ~x01 & ~x02 & ~x03) | (x02 & x03 & x00 & x01)));
  assign z06 = (~x13 & ((x02 & (x00 ? (~x01 & ~x07 & (x04 ? ((~x10 & ((~x12 & ((x09 & ((x03 & x08 & (x14 | x15)) | (~x14 & x15 & ~x16 & ~x03 & ~x08 & x11))) | (~x15 & x16 & ~x11 & ~x14 & ~x08 & ~x09 & ~x03 & x06))) | (x03 & ~x08 & x09 & x15 & ~x16 & ~x11 & ~x14))) | (~x14 & x15 & ~x16 & x11 & x12 & ~x09 & x10 & ~x03 & ~x08)) : (x09 & ~x10 & ((x08 & (x14 | x15) & (x03 | (~x03 & ~x11 & ~x12))) | (~x14 & x15 & ~x16 & x03 & ~x08))))) : ((~x14 & ((~x15 & ((~x06 & ((x01 & ((x03 & ~x04 & ((~x12 & x16 & ~x10 & ~x11 & ~x07 & ~x08 & ~x09) | (~x05 & x07 & ~x16))) | (~x09 & ~x10 & ~x11 & ~x12 & x16 & ~x07 & ~x08 & ~x03 & x04))) | (~x01 & ~x03 & x04 & ~x05 & ~x16))) | (~x01 & ((x05 & x06 & x07 & (x03 ? (x04 | (~x04 & ~x16)) : (x04 & ~x16))) | (~x03 & ~x04 & x16))))) | (~x01 & x03 & ~x04 & ~x07 & x15 & ~x16 & (x08 | (x09 & ~x11 & x12))))) | ((x14 | x15) & (x01 ? (~x03 | (x03 & x04 & ~x06)) : (x03 & ~x04 & ~x07 & ~x10 & ((x09 & (~x08 | (x11 & x12))) | (x08 & ~x11 & ~x12)))))))) | (~x07 & ((x09 & (((x14 | x15) & ((~x02 & ((x00 & ~x01 & ~x10 & ((x03 & x08 & ~x11 & ~x12) | (x04 & ~x08))) | (~x00 & x01 & x03 & ~x11 & ~x12 & ~x08 & x10))) | (~x11 & ~x12 & ~x08 & x10 & ~x03 & ~x04 & ~x00 & x01))) | (~x03 & x04 & x00 & ~x02 & ~x14 & x15 & ~x16 & ~x08 & ~x10))) | (~x02 & x04 & ~x09 & ~x10 & ((x16 & ((~x08 & ~x11 & ~x12 & ~x14 & ~x15 & ((x00 & x06 & (x01 | x03)) | (~x00 & x01 & x03 & ~x06))) | (x00 & ~x01 & ~x03 & x08 & x15))) | (x00 & ~x01 & ~x03 & x08 & x14))))) | (~x00 & ~x14 & ~x15 & x16 & ((~x01 & x03 & x04) | (~x03 & ~x04 & x01 & ~x02))))) | (x07 & ((x13 & ((x02 & (x00 ? (~x01 & x05 & x06 & (x03 ^ x04)) : (x01 & x03 & ~x04 & ~x05 & (x14 ^ x15)))) | (~x00 & x01 & ~x02 & ~x05 & ((~x14 & x15 & ~x16 & ~x03 & ~x04) | (x08 & ((~x03 & ~x04 & (x14 ? ~x15 : (x15 & x16))) | (x03 & x04 & x14 & ~x15))))))) | (x02 & ~x03 & ~x00 & x01 & ~x04 & ~x05 & x08 & x14 & ~x15))) | (x00 & x01 & x02 & x03 & x04);
  assign z07 = (~x01 & ((x07 & x13 & x05 & x06 & ~x03 & ~x04 & x00 & x02) | (x03 & x04 & ~x00 & ~x02 & ~x15 & x16 & ~x13 & ~x14))) | (~x00 & x01 & x02 & ~x04 & (x03 ? (~x05 & x07 & x13 & (x14 ^ x15)) : (~x13 & (x14 | x15 | (~x08 & ~x09 & ~x06 & ~x07 & ~x12 & x16 & ~x10 & ~x11)))));
  assign z08 = (~x01 & ((x07 & x13 & x05 & x06 & ~x03 & ~x04 & x00 & x02) | (x03 & x04 & ~x00 & ~x02 & ~x15 & x16 & ~x13 & ~x14))) | (~x00 & x01 & x02 & ~x04 & (x03 ? (~x05 & x07 & x13 & (x14 ^ x15)) : (~x13 & (x14 | x15 | (~x08 & ~x09 & ~x06 & ~x07 & ~x12 & x16 & ~x10 & ~x11)))));
  assign z09 = (x02 & ((~x13 & ((~x07 & ~x10 & ((~x11 & ((x00 & ~x01 & x09 & ((x03 & x04 & ~x08 & ~x14 & x15 & ~x16) | (~x03 & ~x04 & x08 & ~x12 & (x14 | x15)))) | (~x03 & ~x04 & ~x00 & x01 & ~x06 & ~x08 & ~x09 & ~x12 & x16))) | (x00 & ~x01 & x03 & x04 & x08 & x09 & x11 & ~x12 & (x14 | x15)))) | (~x00 & x01 & ~x03 & ~x04 & (x14 | x15)))) | (x07 & x13 & x05 & x06 & ~x03 & ~x04 & x00 & ~x01))) | (~x15 & x16 & ~x13 & ~x14 & x03 & x04 & ~x00 & ~x01);
  assign z10 = x01 ? ((~x00 & ~x03 & ((~x09 & ~x10 & ((~x02 & x04 & ~x05 & x07 & x08 & x13 & x14 & ~x15 & ~x16 & (x11 ^ x12)) | (~x06 & ~x07 & x02 & ~x04 & ~x08 & ~x11 & ~x12 & ~x13 & x16))) | (x02 & ~x04 & ~x13 & (x14 | x15)))) | (x00 & ~x02 & ~x04 & ~x08 & ~x09 & x06 & ~x07 & ~x10 & ~x11 & ~x12 & ~x15 & x16 & ~x13 & ~x14)) : ((x04 & ((~x13 & ((~x07 & ~x08 & ((x15 & ((~x14 & ~x16 & ((x00 & x02 & ~x03 & x11 & (x09 ? (~x10 & ~x12) : (x10 & x12))) | (x09 & ~x10 & ~x02 & x03))) | (~x00 & ~x02 & x03 & x09 & ~x10))) | (~x00 & ~x02 & x03 & x09 & ~x10 & x14))) | (~x00 & x03 & ~x14 & ~x15 & x16))) | (~x00 & ~x02 & x03 & ~x05 & x07 & x08 & ~x09 & ~x10 & x13 & (x11 ^ x12) & (x14 ? ~x15 : (x15 & x16))))) | (x00 & ~x04 & ((x06 & ((x02 & ((~x03 & x05 & x07 & x13) | (~x07 & ~x08 & ~x09 & ~x10 & ~x11 & ~x14 & ~x15 & x16 & ~x12 & ~x13))) | (~x14 & ~x15 & x16 & ~x11 & ~x12 & ~x13 & ~x08 & ~x09 & ~x10 & ~x02 & x03 & ~x07))) | (~x02 & ~x07 & ~x08 & x09 & ~x10 & ~x13 & (x14 | x15)))));
  assign z11 = x04 ? ((~x13 & ((~x07 & ((~x10 & ((~x08 & ((~x02 & ((~x14 & ((~x09 & ~x11 & ~x12 & ~x15 & ((x16 & ((x00 & x06 & (x01 | x03)) | (~x00 & x01 & x03 & ~x06))) | (~x05 & ~x06 & ~x16 & ~x00 & x01 & x03))) | (x00 & ~x03 & x09 & x15 & ~x16))) | (x00 & ~x01 & x09 & (x14 | x15)))) | (~x01 & x02 & ~x03 & (x00 ? (~x12 & ~x14 & ((x06 & ~x09 & ~x11 & ~x15 & x16) | (x15 & ~x16 & x09 & x11))) : (x09 & (x14 | x15)))))) | (~x01 & x08 & ((x02 & ~x11 & ~x12 & (x00 ? (x03 & x09 & (x14 | x15)) : (~x03 & ~x09 & (x14 | x16)))) | (x00 & ~x02 & ~x03 & ~x09 & (x14 | (x15 & x16))))))) | (~x00 & ~x02 & x03 & (((x14 | x15) & ((~x01 & x08) | (x10 & ~x11 & ~x12 & x01 & ~x08 & x09))) | (~x01 & ~x08 & x09 & x10 & ~x14 & x15 & ~x16 & ~x11 & x12))) | (~x14 & x15 & ~x16 & x10 & x11 & x12 & x00 & ~x01 & x02 & ~x03 & ~x08 & ~x09))) | (~x00 & ~x14 & ~x15 & ((~x02 & ((x06 & x07 & x08 & ~x01 & x03 & x05) | (x01 & ~x03 & x16))) | (~x01 & ((x03 & (x16 | (x06 & x07 & x02 & x05))) | (x02 & ~x03 & (x16 | (x07 & ~x16 & x05 & x06))))))))) | (x02 & x03 & x00 & x01) | (x07 & x13 & ((~x05 & ((~x14 & x15 & ((~x09 & ((~x10 & (x00 ? (x01 & x02 & ~x03 & ((~x12 & x16 & x08 & ~x11) | (x11 & x12 & ~x16))) : (~x01 & ~x02 & x03 & x08 & x16 & (~x12 | (~x11 & x12))))) | (x10 & ~x11 & ~x12 & ~x16 & x02 & ~x03 & x00 & x01))) | (x02 & ((~x00 & ((x01 & ~x03) | (~x01 & x03 & x08 & x16))) | (x00 & x01 & ~x03 & ~x08 & ~x16))))) | (x02 & x14 & ~x15 & ((x01 & ~x03 & (~x00 | (x00 & x08 & ~x09 & ~x10 & x16 & (x11 ^ x12)))) | (x03 & x08 & ~x00 & ~x01))))) | (x00 & ~x01 & x02 & x03 & x05 & x06)))) : ((~x13 & ((~x07 & ((~x10 & ((~x08 & ((~x09 & ~x11 & ~x12 & ((~x14 & ~x15 & ((x00 & x06 & x16 & (x01 ? (~x02 & x03) : ~x03)) | (~x00 & x01 & ~x02 & ~x06 & ~x16 & ~x03 & ~x05))) | (~x00 & x01 & x02 & ~x03 & ~x06 & x16))) | (x00 & ~x01 & ~x02 & x03 & x09 & (x14 | x15)))) | (x00 & ~x02 & x08 & (x01 ? (x03 & x09 & (x14 | x15)) : (~x03 & ~x09 & ~x11 & (x14 | (x15 & x16))))))) | (~x00 & x01 & ~x03 & ~x08 & x09 & x10 & ~x11 & ~x12 & (x14 | x15)))) | (~x00 & x02 & ((x01 & ~x03 & (x14 | x15)) | (~x15 & ~x16 & ~x06 & ~x14 & ~x01 & x03 & ~x05))) | (~x14 & ~x15 & ~x16 & ~x06 & x07 & x00 & ~x01 & ~x02 & ~x03 & ~x05))) | (~x03 & x07 & ((~x00 & x01 & ~x05 & ((x14 & ~x15 & x02 & x08) | (~x14 & x15 & ~x16 & ~x02 & x13))) | (x00 & ~x01 & x02 & x05 & x06 & x13))));
  assign z12 = (~x00 & ((x04 & (x01 ? ((~x03 & ~x05 & x07 & x13 & (x02 ? (x14 ^ x15) : (x08 & ~x09 & ~x10 & x14 & ~x15 & ~x16 & (x11 ^ x12)))) | (~x10 & ~x11 & ~x12 & ~x15 & x16 & ~x13 & ~x14 & ~x07 & ~x08 & ~x09 & ~x02 & x03 & ~x06)) : ((~x13 & ((~x14 & ((~x15 & ((x03 & (x16 | (~x02 & ~x16 & ((~x05 & ~x06) | (x05 & x06 & x07 & ~x08))))) | (x06 & x07 & ~x16 & x02 & ~x03 & x05))) | (~x02 & x03 & ~x07 & ~x08 & x09 & x10 & ~x11 & x12 & x15 & ~x16))) | (~x02 & x03 & ~x07 & ~x08 & x09 & ~x10 & (x14 | x15)))) | (~x02 & x03 & ~x05 & x07 & x08 & ~x09 & ~x10 & x13 & x16 & ((~x11 & x12 & (x14 ^ x15)) | (~x12 & ((~x14 & x15) | (x11 & x14 & ~x15)))))))) | (~x14 & ((x01 & ~x04 & ~x05 & x07 & ~x16 & ((~x02 & ~x03 & x13 & x15) | (x02 & x03 & ~x06 & ~x13 & ~x15))) | (~x13 & ~x15 & x16 & ~x01 & ~x02 & x03))) | (x01 & ~x03 & ~x04 & ~x13 & (((x14 | x15) & (x02 | (x10 & ~x11 & ~x12 & ~x07 & ~x08 & x09))) | (~x09 & ~x10 & ~x11 & ~x12 & x16 & ~x07 & ~x08 & x02 & ~x06))))) | (x00 & ((x06 & ((~x01 & x02 & ~x03 & x05 & x07 & x13) | (~x14 & ~x15 & x16 & ~x11 & ~x12 & ~x13 & ~x08 & ~x09 & ~x10 & ~x02 & ~x04 & ~x07))) | (~x01 & ~x07 & ~x13 & ((x02 & ~x03 & x04 & ~x08 & ~x09 & ~x14 & x15 & ~x16 & x10 & x11 & x12) | (x09 & ~x10 & (((x14 | x15) & ((~x02 & ~x03 & ~x04 & ~x08) | (x02 & x03 & x04 & x08 & x11 & ~x12))) | (~x14 & x15 & ~x16 & x11 & ~x12 & x04 & ~x08 & x02 & ~x03))))) | (x03 & x04 & x01 & x02))) | (~x01 & ~x02 & x03 & x04 & ~x07 & ~x08 & ~x14 & x15 & ~x16 & x09 & ~x10 & ~x13);
  assign z13 = (~x01 & ((~x13 & ((x03 & (x00 ? (~x07 & x09 & ~x10 & (x14 | x15) & ((~x02 & ~x04 & (~x08 | (x08 & ~x11 & ~x12))) | (x02 & x04 & x08 & ~x11 & ~x12))) : ((~x14 & ((~x15 & ((x02 & ((x06 & x07 & x04 & x05) | (~x06 & ~x16 & ~x04 & ~x05))) | x16 | (~x02 & x04 & ~x16 & ((~x05 & ~x06) | (x05 & x06 & x07 & ~x08))))) | (x02 & ~x04 & ~x07 & x15 & ~x16 & (x08 | (x09 & ~x11 & x12))))) | (~x07 & (((x14 | x15) & ((x08 & ((~x02 & x04) | (~x10 & ~x11 & ~x12 & x02 & ~x04))) | (x02 & ~x04 & x09 & ((~x08 & (~x10 | (x10 & ~x11 & ~x12))) | (~x10 & x11 & x12))))) | (x02 & ~x04 & x08 & ~x09 & ~x10 & ~x11 & x12 & (x14 | (x15 & x16)))))))) | (~x03 & ((~x07 & ((~x10 & ((~x09 & ((x08 & ((x04 & (x00 ? (~x02 & (x14 | (x15 & x16))) : (x02 & ~x11 & ~x12 & (x14 | x16)))) | (x00 & ~x02 & ~x04 & ~x11 & (x14 | (x15 & x16))))) | (x00 & x06 & ~x08 & ~x11 & ~x12 & ~x14 & ~x15 & x16 & (~x04 | (x02 & x04))))) | (x02 & x04 & ~x08 & x09 & ((~x00 & (x14 | x15)) | (~x14 & x15 & ~x16 & x00 & x11 & ~x12))))) | (~x14 & x15 & ~x16 & x10 & x11 & x12 & x04 & ~x08 & ~x09 & x00 & x02))) | (~x14 & ~x15 & ((x04 & x16 & ~x00 & x02) | (x07 & ~x16 & ~x05 & ~x06 & x00 & ~x02 & ~x04))))) | (x00 & ~x02 & x04 & ~x07 & ~x08 & x09 & ~x10 & (x14 | x15)))) | (x07 & x13 & ((x02 & (x00 ? (x05 & x06 & (x04 | (~x03 & ~x04))) : (x03 & x04 & ~x05 & x08 & (x14 ? ~x15 : (x15 & x16))))) | (~x00 & ~x02 & x03 & x04 & ~x05 & x08 & ~x09 & ~x10 & x14 & ~x15 & x16 & (x11 ^ x12)))) | (~x03 & ~x04 & ~x00 & ~x02))) | (x04 & ((~x09 & ((~x10 & ((~x15 & ((x01 & ((~x05 & ((~x03 & x07 & x08 & x13 & x14 & (x11 ^ x12) & (x00 ? (x02 & x16) : (~x02 & ~x16))) | (~x00 & ~x02 & x03 & ~x06 & ~x07 & ~x08 & ~x11 & ~x12 & ~x13 & ~x14 & ~x16))) | (~x02 & ~x07 & ~x08 & ~x11 & ~x12 & ~x13 & ~x14 & x16 & (x00 ? x06 : (x03 & ~x06))))) | (x00 & ~x02 & x03 & x06 & ~x07 & ~x08 & ~x11 & ~x12 & ~x13 & ~x14 & x16))) | (x00 & x01 & x02 & ~x03 & ~x05 & x07 & x13 & ~x14 & x15 & ((~x12 & x16 & x08 & ~x11) | (x11 & x12 & ~x16))))) | (x00 & x01 & x02 & ~x03 & ~x05 & x07 & x10 & ~x11 & ~x12 & x15 & ~x16 & x13 & ~x14))) | (~x08 & ((x15 & ((x00 & ~x03 & ~x14 & ~x16 & ((x01 & x02 & ~x05 & x07 & x13) | (x09 & ~x10 & ~x13 & ~x02 & ~x07))) | (~x00 & x01 & ~x02 & x03 & ~x07 & ~x11 & ~x12 & ~x13 & x09 & x10))) | (~x00 & x01 & ~x02 & x03 & ~x07 & x09 & x10 & ~x11 & ~x12 & ~x13 & x14))) | (~x15 & x16 & ~x13 & ~x14 & ~x02 & ~x03 & ~x00 & x01))) | (~x04 & ((x01 & ((~x13 & (((x14 | x15) & ((~x00 & x02 & ~x03) | (x00 & ~x02 & x03 & x09 & ~x10 & ~x07 & x08))) | (~x14 & ~x15 & ~x16 & ~x06 & x07 & x03 & ~x05 & ~x00 & x02))) | (x02 & ((x00 & x03) | (~x00 & ~x03 & ~x05 & x14 & ~x15 & x07 & x08))))) | (~x10 & ~x11 & ~x12 & ~x15 & x16 & ~x13 & ~x14 & ~x08 & ~x09 & x06 & ~x07 & x00 & ~x02 & ~x03)));
  assign z14 = (~x13 & ((~x01 & ((~x00 & (x02 ? ((~x04 & ((~x16 & (x03 ? (~x07 & ~x14 & x15 & (x08 | (x09 & ~x11 & x12))) : (x05 ? (x06 & x07) : ~x06))) | (x03 & ~x07 & ((~x08 & x09 & x10 & ~x11 & ~x12 & (x14 | x15)) | (~x10 & (((x14 | x15) & ((x09 & (~x08 | (x11 & x12))) | (x08 & ~x11 & ~x12))) | (x08 & ~x09 & ~x11 & x12 & (x14 | (x15 & x16))))))))) | (~x15 & x16 & x03 & ~x14)) : (x04 & ((~x08 & ((x03 & ~x14 & ~x16 & ((~x07 & x09 & x10 & ~x11 & x12 & x15) | (x05 & x06 & x07 & ~x15))) | (~x07 & x09 & ~x10 & x11 & (x14 | x15)))) | (~x14 & ~x15 & ~x16 & x03 & ~x05 & ~x06))))) | (~x07 & ((x00 & ((x02 & ~x03 & x04 & ~x08 & ~x09 & ~x14 & x15 & ~x16 & x10 & x11 & x12) | (~x10 & ((x09 & ((x15 & (x02 ? ((x03 & ~x04 & x08) | (~x03 & x04 & ~x08 & x11 & ~x12 & ~x14 & ~x16)) : ((x03 & ((~x11 & ~x12 & ~x04 & x08) | (~x14 & ~x16 & ~x08 & x11))) | (~x04 & ~x08 & x11) | (~x03 & x04 & x08 & ~x11 & ~x12)))) | (x14 & ((~x04 & (x02 ? (x03 & x08) : ((x03 & x08 & ~x11 & ~x12) | (~x08 & x11)))) | (x08 & ~x11 & ~x12 & ~x02 & ~x03 & x04))))) | (x06 & ~x08 & ~x09 & ~x11 & ~x12 & ~x14 & ~x15 & x16 & ((~x03 & ~x04) | (~x02 & (x03 ^ x04)))))))) | (x02 & x03 & x04 & x06 & ~x08 & ~x09 & ~x14 & ~x15 & x16 & ~x10 & ~x11 & ~x12))))) | (~x04 & (((x14 | x15) & ((~x00 & ~x03 & (x02 | (x01 & ~x07 & ~x08 & ~x11 & ~x12 & x09 & x10))) | (x09 & ~x10 & ~x07 & x08 & x00 & x01 & ~x02 & x03))) | (~x00 & x01 & x02 & ~x03 & ~x06 & ~x07 & ~x11 & ~x12 & x16 & ~x08 & ~x09 & ~x10))) | (~x00 & x01 & x04 & ~x06 & ~x14 & ~x15 & ((~x02 & ~x07 & ~x08 & ~x09 & ~x10 & ~x11 & ~x12 & (x03 ? x16 : (~x05 & ~x16))) | (x02 & ~x03 & ~x05 & x07 & ~x16))))) | (~x00 & ((~x05 & x07 & x08 & ((~x03 & ((~x04 & (x14 ? ~x15 : (x15 & x16)) & (x01 ? (~x02 & x13) : x02)) | (x01 & ~x02 & x04 & ~x09 & ~x10 & x14 & ~x15 & ~x16 & x11 & ~x12 & x13))) | (~x02 & x03 & x13 & ((~x01 & x04 & ~x09 & ~x10 & ~x12 & ((~x14 & x15 & x16) | (x11 & x14 & ~x15))) | (x14 & ~x15 & ~x16 & x01 & ~x04))))) | (~x01 & ~x02 & ~x03))) | (x00 & x01 & x02 & x03 & ~x04);
endmodule