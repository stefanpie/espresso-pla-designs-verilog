module pla__apex2 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38,
    z0, z1, z2  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38;
  output z0, z1, z2;
  assign z0 = ~x28 & ((~x23 & ((~x16 & ~x27 & (((~x13 | ~x14) & (((~x12 | ~x17) & (((x34 ? ~x24 : x35) & ((x07 & ~x09 & x31 & (x21 | ~x29)) | (~x07 & ~x29 & ~x30 & x36 & (~x08 | ~x32)) | (x29 & (x22 | (x20 & ~x21))))) | (~x24 & ((~x26 & ((~x29 & ~x30 & x36 & ((~x07 & (~x08 | ~x32)) | (~x08 & ~x31 & ~x35))) | (x29 & (x22 | (~x21 & (x00 | (x20 & ~x22))))) | (x07 & ~x09 & x31))) | (~x08 & ~x29 & ~x30 & ~x31 & x34 & ~x35 & x36))))) | (x36 & (~x08 | ~x32) & ((~x24 & (~x07 | (~x31 & ~x35)) & ((~x26 & ((~x02 & ((~x04 & ~x05 & ~x06 & ((~x01 & ~x17 & (~x21 | ~x29)) | (~x12 & ~x29))) | (~x17 & ~x21 & ~x30))) | (~x12 & ~x21 & (~x30 | (~x04 & ~x05 & ~x06 & x29))))) | (~x02 & ~x04 & ~x05 & ~x06 & ~x29 & x34 & (~x12 | (~x01 & ~x17))))) | (~x02 & ~x04 & ~x05 & ~x06 & ~x07 & ~x29 & ~x34 & x35 & (~x12 | (~x01 & ~x17))))) | (x02 & ~x12 & ~x20 & ~x21 & ~x24 & ~x26 & x29))) | (~x17 & ((~x09 & (x13 ? ~x14 : (~x10 | (x03 & ~x18) | (~x11 & ~x19))) & ((~x04 & ~x05 & ~x06 & x36 & (~x08 | ~x32) & ((~x24 & ((((~x21 & ~x26 & x29) | (~x02 & ~x29 & x34)) & (~x07 | ~x35)) | (~x02 & ~x26 & ~x29 & ~x35))) | (~x02 & ~x07 & ~x29 & ~x34 & x35))) | (x02 & ~x21 & ~x24 & ~x26 & x29))) | ((x34 ? ~x24 : x35) & (x21 | ~x29) & ((~x14 & ((x07 & x10 & x13 & x31) | (x25 & x33))) | (~x13 & ((x07 & x10 & x31 & ((x03 & ~x18) | (~x11 & ~x19))) | (x14 & x33))))) | (~x24 & ~x26 & ((~x14 & ((x07 & x10 & x13 & x31) | (x25 & x33))) | (~x13 & ((x07 & x10 & x31 & ((x03 & ~x18) | (~x11 & ~x19))) | (x14 & x33))))))) | (~x12 & (((x34 ? ~x24 : x35) & (x21 | ~x29) & ((~x14 & ((x07 & x10 & x13 & x31) | (x25 & x33))) | (~x13 & ((x07 & x10 & x31 & ((x03 & ~x18) | (~x11 & ~x19))) | (x14 & x33))))) | (~x24 & ~x26 & ((~x14 & ((x07 & x10 & x13 & x31) | (x25 & x33))) | (~x13 & ((x07 & x10 & x31 & ((x03 & ~x18) | (~x11 & ~x19))) | (x14 & x33))))))))) | (~x24 & ~x30 & ~x31 & ~x32 & x34 & ((x33 & (x21 | ~x29) & (x14 | x25)) | (x29 & (x22 | (x20 & ~x21))) | (~x29 & x36 & (~x07 | ~x35)))))) | (~x30 & ~x31 & ~x32 & ~x34 & (((x35 | (~x24 & ~x26)) & ((x29 & (x22 | (x20 & ~x21))) | (x33 & (x21 | ~x29) & (x14 | x25)))) | (~x29 & x36 & ((~x07 & x35) | (~x24 & ~x26 & ~x35))))));
  assign z1 = ~x28 & ((~x23 & ((~x16 & ~x27 & (((~x13 | ~x14) & ((~x24 & ((~x26 & ((x29 & ((x02 & ~x20 & (~x17 | (~x12 & ~x21))) | ((~x12 | ~x17) & (x22 | (x21 & ~x22))))) | ((~x12 | ~x17) & ((x25 & x33) | (x07 & x31))))) | (x34 & (~x12 | ~x17) & ((((x25 & x33) | (x07 & x31)) & (x20 | ~x29)) | (x29 & (x21 | x22)))))) | (~x34 & x35 & (~x12 | ~x17) & ((((x25 & x33) | (x07 & x31)) & (x20 | ~x29)) | (x29 & (x21 | x22)))))) | (x37 & (((~x08 | ~x32) & ((~x24 & (((~x07 | ~x35) & ((~x04 & ~x05 & ~x06 & ((~x02 & ~x29 & x34) | (~x26 & x29 & ~x00 & ~x20)) & (((~x14 | (~x13 & ~x33)) & (~x12 | (~x17 & (~x01 | (~x09 & (~x10 | (x03 & ~x18) | (~x11 & ~x19))))))) | (~x09 & x13 & ~x14 & ~x17))) | (~x00 & ~x20 & ~x26 & ~x30 & (~x12 | ~x17) & (~x14 | (~x13 & ~x33))))) | (~x02 & ~x04 & ~x05 & ~x06 & ~x26 & ~x29 & ~x35 & (((~x14 | (~x13 & ~x33)) & (~x12 | (~x17 & (~x01 | (~x09 & (~x10 | (x03 & ~x18) | (~x11 & ~x19))))))) | (~x09 & x13 & ~x14 & ~x17))))) | (~x02 & ~x04 & ~x05 & ~x06 & ~x07 & ~x29 & ~x34 & x35 & (((~x14 | (~x13 & ~x33)) & (~x12 | (~x17 & (~x01 | (~x09 & (~x10 | (x03 & ~x18) | (~x11 & ~x19))))))) | (~x09 & x13 & ~x14 & ~x17))))) | (~x29 & ~x30 & (((x34 ? ~x24 : x35) & (~x14 | (~x13 & ~x33)) & (~x12 | ~x17) & ((~x07 & ~x08) | (x31 & ~x32))) | (~x24 & (~x14 | (~x13 & ~x33)) & (~x12 | ~x17) & ((~x08 & ~x35 & (~x26 | x34)) | (~x26 & x31 & ~x32))))))))) | (~x24 & ~x30 & ~x31 & ~x32 & x34 & ((~x29 & ((x25 & x33) | (x37 & (~x07 | ~x35) & (~x14 | ~x33)))) | (x29 & (x21 | x22)) | (x20 & x25 & x33))))) | (~x30 & ~x31 & ~x32 & ~x34 & ((~x29 & ((x37 & (~x14 | ~x33) & ((~x07 & x35) | (~x24 & ~x26 & ~x35))) | (x25 & x33 & (x35 | (~x24 & ~x26))))) | ((x35 | (~x24 & ~x26)) & ((x29 & (x21 | x22)) | (x20 & x25 & x33))))));
  assign z2 = ~x28 & ((~x24 & ((~x26 & ((~x22 & ((x29 & ((~x16 & ~x23 & ~x27 & (x21 | (x20 & ~x21)) & (~x13 | ~x14) & (~x12 | ~x17)) | x16 | (x13 & x14) | (x12 & x17) | x23 | x27)) | (x38 & (~x25 | ~x33) & (~x08 | ~x32) & (((~x07 | (~x31 & ~x35)) & ((~x30 & (~x02 | (x12 & (x09 | (x10 & ~x13 & (~x03 | x18) & (x11 | x19)))))) | (~x02 & ~x04 & ~x05 & ~x06 & ((~x09 & ((x03 & ~x18) | (~x11 & ~x19) | ~x10 | x13)) | ~x01 | ~x12)))) | (x09 & ~x35 & ((~x02 & (~x30 | (~x04 & ~x05 & ~x06 & (~x01 | ~x12)))) | (x12 & ~x30)) & (~x10 | (~x13 & (~x03 | x18) & (x11 | x19)))))))) | ((x16 | (x13 & x14) | (x12 & x17) | x23 | x27) & (x30 | x31 | x32)) | (x14 & x33) | (~x29 & x38 & (~x25 | ~x33) & (~x08 | ~x32) & (((~x07 | (~x31 & ~x35)) & (~x30 | (~x02 & ~x04 & ~x05 & ~x06 & ((~x09 & ((x03 & ~x18) | (~x11 & ~x19) | ~x10 | x13)) | ~x01 | ~x12)))) | (x09 & ~x35 & (~x10 | (~x13 & (~x03 | x18) & (x11 | x19))) & (~x30 | (~x02 & ~x04 & ~x05 & ~x06 & (~x01 | ~x12)))))))) | (x34 & ((~x29 & ((~x13 & ((x14 & ~x16 & ~x23 & ~x27 & x33 & (~x12 | ~x17)) | (x09 & ~x35 & x38 & (~x25 | ~x33) & (x11 | x19) & (~x08 | ~x32) & (~x03 | x18) & (~x30 | (~x02 & ~x04 & ~x05 & ~x06 & (~x01 | ~x12)))))) | ((x30 | x31 | x32) & (x16 | (x13 & x14) | x27 | (x12 & x17))) | (x38 & (~x25 | ~x33) & (~x08 | ~x32) & (((~x07 | (~x31 & ~x35)) & (~x30 | (~x02 & ~x04 & ~x05 & ~x06 & ((~x09 & ((x03 & ~x18) | (~x11 & ~x19) | ~x10 | x13)) | ~x01 | ~x12)))) | (x09 & ~x10 & ~x35 & (~x30 | (~x02 & ~x04 & ~x05 & ~x06 & (~x01 | ~x12)))))) | x23 | (x14 & ~x23 & ~x30 & ~x31 & ~x32 & x33))) | (~x22 & x29 & (x20 | x21)) | (x22 & (((x30 | x31 | x32) & (x16 | (x13 & x14) | x27 | (x12 & x17))) | x23 | (x14 & x33))))))) | (~x34 & x35 & ((~x29 & ((x14 & ((x33 & ((~x30 & ~x31 & ~x32) | (~x13 & ~x16 & ~x23 & ~x27 & (~x12 | ~x17)))) | (x13 & (x30 | x31 | x32)))) | ((x30 | x31 | x32) & (x23 | x27 | x16 | (x12 & x17))) | (~x07 & x38 & (~x25 | ~x33) & (~x08 | ~x32) & (~x30 | (~x02 & ~x04 & ~x05 & ~x06 & ((~x09 & ((x03 & ~x18) | (~x11 & ~x19) | ~x10 | x13)) | ~x01 | ~x12)))))) | (~x22 & x29 & (x20 | x21)) | (x22 & ((x14 & x33) | ((x16 | (x13 & x14) | (x12 & x17) | x23 | x27) & (x30 | x31 | x32)))))));
endmodule