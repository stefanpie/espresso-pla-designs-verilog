module pla__xparc ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71, z72  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71, z72;
  assign z00 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & (x00 ? (~x01 & ~x02 & ~x14 & ((~x12 & x13 & ((x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17)) & (x03 ? (~x04 & ~x05) : (~x04 | (x04 & ~x05)))) | (~x03 & ~x04 & ~x05 & x15 & ~x18 & x19 & ~x16 & ~x17))) | (~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19))) : ((x13 & ((x15 & ((~x17 & ((~x02 & ((~x12 & ~x14 & ~x18 & (((~x01 | (x01 & x16 & ~x19)) & (x05 ? ~x03 : x04)) | (~x03 & ~x04 & ((x01 & (x19 | (~x05 & ~x19))) | (~x01 & ~x05 & ~x16 & x40))) | (x01 & x04 & ~x16 & x19))) | (~x01 & ~x03 & ~x04 & ~x05 & x12 & x14 & x40 & (x16 | (~x16 & x19))))) | (~x12 & ~x14 & ~x18 & (((~x01 | (x01 & x16 & ~x19)) & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))))) | (x01 & ~x16 & x19 & ((x02 & (~x03 | (x03 & x04))) | (x03 & ~x04))))))) | (~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x14 & x40 & (x12 | (~x12 & ~x16 & x17 & x18 & x19))))) | (~x15 & ((~x01 & ((~x14 & ((~x12 & x16 & x17 & x18 & x19 & ((x03 & (~x04 | (x04 & x05))) | (~x02 & ((x04 & ~x05) | (~x03 & (x05 | (~x04 & ~x05 & x40))))))) | (~x02 & ~x03 & ~x04 & ~x05 & x12 & x40 & ((x24 & x25 & x28) | (~x28 & ~x31))))) | (~x02 & ~x03 & ~x04 & ~x05 & x12 & x14 & x40 & ((x18 & x19 & ~x16 & x17) | (~x17 & ~x18 & ~x19))))) | (~x12 & ~x14 & x16 & x17 & x18 & x19 & (x02 ? (~x03 | (x03 & ((x04 & ~x05) | (x01 & (~x04 | (x04 & x05)))))) : x01)))) | (~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x12 & ~x14 & x16 & ~x17 & ~x18 & x40))) | (~x01 & ~x02 & ~x04 & x12 & ~x13 & ((~x03 & ((~x05 & x40 & (x14 | (~x14 & ((~x16 & (x15 ? (x19 ? ~x18 : x17) : (~x18 & ~x19))) | (~x15 & x17 & ((x18 & x19) | (x16 & (x18 ^ x19)))))))) | (x05 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ~x19))) | (~x16 & x17 & ~x18 & ~x19 & ~x14 & ~x15 & x03 & ~x05)))));
  assign z02 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x36 & x40 & (x13 ? (x14 ? (~x16 & ((x15 & ~x17) | (~x18 & x19 & ~x15 & x17))) : (~x15 & ~x28)) : x14);
  assign z03 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x36 & x40 & ((x14 & (~x13 | (~x16 & ~x17 & x13 & x15))) | (x13 & ~x14 & ~x15 & (~x28 | (x28 & (~x24 | (x24 & ~x25))))));
  assign z04 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x14 & (x00 ? (~x01 & ~x02 & ((~x12 & x13 & ((x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17)) & (x03 ? (~x04 & ~x05) : (~x04 | (x04 & ~x05)))) | (~x03 & ~x04 & ~x05 & x15 & ~x18 & x19 & ~x16 & ~x17))) | (~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19))) : ((~x02 & ((~x01 & (x05 ? (~x12 & x13 & ((x15 & ~x17 & ~x18 & ((~x03 & (~x16 ^ x19)) | (x04 & (~x16 ^ ~x19)))) | (x17 & x18 & x19 & x04 & ~x15 & x16))) : ((x13 & ((~x12 & ((~x17 & ~x18 & ((x15 & ((x04 & (~x16 ^ x19)) | (~x03 & ~x04 & ~x16 & x19 & x40))) | (~x03 & ~x04 & x16 & x40 & (~x19 | (~x15 & x19))))) | (~x03 & ~x04 & x17 & x18 & x19 & x40 & (x15 ^ x16)))) | (~x03 & ~x04 & x12 & x40 & ((~x15 & x24 & x25 & x27 & x28) | (x15 & x29))))) | (~x04 & x12 & ~x13 & x17 & ~x19 & ((~x03 & x40 & (x15 ? (~x16 & x18) : (~x16 ^ x18))) | (~x16 & ~x18 & x03 & ~x15)))))) | (~x12 & x13 & ((x15 & ~x17 & ~x18 & ((x01 & ((x05 & (x03 ? (x04 & (~x16 ^ ~x19)) : (x16 & ~x19))) | (~x03 & ~x04 & (x19 | (~x05 & ~x19))))) | (x03 & x04 & ~x05 & (~x16 ^ ~x19)))) | (x17 & x18 & x19 & x01 & ~x15 & x16))))) | (~x12 & x13 & (x15 ? (~x17 & ~x18 & ((x04 & ((x03 & ((x02 & ((~x01 & ~x05) | ((~x16 ^ ~x19) & (x05 | (x01 & ~x05))))) | (~x01 & x05 & (~x16 ^ x19)))) | (x01 & ~x03 & (x16 ? (~x19 & (~x05 | (x02 & x05))) : x19)))) | (~x01 & (x03 ? ~x04 : x02)) | (x01 & ~x04 & (~x16 ^ ~x19) & (x03 | (x02 & ~x03))))) : (x16 & x17 & x18 & x19 & (x03 ? (((~x04 | (x04 & ~x05)) & (~x01 | (x01 & x02))) | (x02 & x04 & x05)) : x02))))))) | (~x03 & ~x04 & ~x05 & ~x00 & ~x01 & ~x02 & x12 & x13 & x14 & x15 & ~x16 & ~x17 & x40));
  assign z05 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x03 & ~x04 & ~x05 & ~x00 & ~x01 & ~x02 & x12 & x13 & x14 & x15 & ~x16 & ~x17 & x40) | (~x14 & ((x13 & (x00 ? (~x01 & ~x02 & ~x12 & ((x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17)) & (x03 ? (~x04 & ~x05) : (~x04 | (x04 & ~x05)))) | (~x03 & ~x04 & ~x05 & x15 & ~x18 & x19 & ~x16 & ~x17))) : ((~x02 & ((~x01 & ((~x03 & ((~x12 & ((~x17 & ~x18 & ((x15 & ((x05 & (~x16 ^ x19)) | (~x04 & ~x05 & ~x16 & x19 & x40))) | (~x04 & ~x05 & x16 & x40 & (~x19 | (~x15 & x19))))) | (~x04 & ~x05 & x17 & x18 & x19 & x40 & (x15 ^ x16)))) | (~x04 & ~x05 & x12 & x40 & (x15 ? x29 : (~x28 | (x28 & (~x24 | (x24 & (~x25 | (x25 & x27)))))))))) | (x04 & ~x12 & ((x15 & ~x17 & ~x18 & (x05 ? (~x16 ^ ~x19) : (~x16 ^ x19))) | (x17 & x18 & x19 & x05 & ~x15 & x16))))) | (~x12 & ((x15 & ~x17 & ~x18 & ((x01 & ((x05 & (x03 ? (x04 & (~x16 ^ ~x19)) : (x16 & ~x19))) | (~x03 & ~x04 & (x19 | (~x05 & ~x19))))) | (x03 & x04 & ~x05 & (~x16 ^ ~x19)))) | (x17 & x18 & x19 & x01 & ~x15 & x16))))) | (~x12 & (x15 ? (~x17 & ~x18 & ((x04 & ((x03 & ((x02 & ((~x01 & ~x05) | ((~x16 ^ ~x19) & (x05 | (x01 & ~x05))))) | (~x01 & x05 & (~x16 ^ x19)))) | (x01 & ~x03 & (x16 ? (~x19 & (~x05 | (x02 & x05))) : x19)))) | (~x01 & (x03 ? ~x04 : x02)) | (x01 & ~x04 & (~x16 ^ ~x19) & (x03 | (x02 & ~x03))))) : (x16 & x17 & x18 & x19 & (x03 ? (((~x04 | (x04 & ~x05)) & (~x01 | (x01 & x02))) | (x02 & x04 & x05)) : x02))))))) | (~x01 & ~x02 & ~x04 & ~x05 & x12 & ~x13 & x17 & ~x19 & ((~x00 & ((~x03 & x40 & (x15 ? (~x16 & x18) : (~x16 ^ x18))) | (~x16 & ~x18 & x03 & ~x15))) | (x00 & ~x03 & ~x15 & ~x16 & ~x18))))));
  assign z06 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x03 & ~x04 & ~x05 & ~x00 & ~x01 & ~x02 & x12 & x13 & x14 & x15 & ~x16 & ~x17 & x40) | (~x14 & ((x13 & (x00 ? (~x01 & ~x02 & ~x03 & ~x12 & ((x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17)) & (~x04 | (x04 & ~x05))) | (~x18 & x19 & ~x16 & ~x17 & ~x04 & ~x05 & x15))) : ((~x01 & ((~x12 & (x15 ? ((~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))) | (~x02 & (x05 ? ~x03 : x04)))) | (~x04 & ~x05 & ~x02 & ~x03 & ~x16 & x17 & x18 & x19 & x40)) : (x16 & ((x17 & x18 & x19 & ((x03 & (~x04 | (x04 & x05))) | (~x02 & (x05 ? ~x03 : x04)))) | (~x02 & ~x03 & ~x04 & ~x18 & x40 & ~x05 & ~x17))))) | (~x02 & ~x03 & ~x04 & ~x05 & x12 & x40 & (x15 ? x29 : (~x28 | (x28 & (~x24 | (x24 & (~x25 | (x25 & x27)))))))))) | (~x12 & ((x01 & ((x16 & (x15 ? (~x17 & ~x18 & ~x19 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))) | (~x02 & (x05 ? ~x03 : x04)))) : (x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))) | (x15 & ~x17 & ~x18 & ((x19 & ((~x02 & ~x03 & ~x04) | (~x16 & ((x02 & (~x03 | (x03 & x04))) | (x03 & ~x04) | (~x02 & x04))))) | (~x02 & ~x03 & ~x04 & ~x05 & ~x19))))) | (x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05)))))))) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & x12 & ~x13 & x17 & ~x19 & ((~x05 & x18 & x40 & (x15 ^ x16)) | (~x16 & ~x18 & x05 & ~x15))))));
  assign z07 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x14 & (x00 ? (~x01 & ~x02 & ~x03 & ((~x12 & x13 & ((x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17)) & (~x04 | (x04 & ~x05))) | (~x18 & x19 & ~x16 & ~x17 & ~x04 & ~x05 & x15))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & ~x04 & ~x05 & x12 & ~x13))) : ((~x01 & ((x13 & ((~x12 & ((~x18 & ((~x17 & ((x15 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))) | (~x02 & ((x04 & ~x05) | (~x03 & (x05 | (~x16 & x40 & ~x04 & ~x05))))))) | (~x02 & ~x03 & ~x04 & ~x05 & x16 & x40))) | (~x02 & ~x03 & ~x04 & ~x15 & x16 & x17 & (x05 ? ~x19 : x40)))) | (~x15 & x16 & x18 & x19 & ((x17 & ((x03 & (~x04 | (x04 & x05))) | (~x02 & (x05 ? ~x03 : x04)))) | (~x04 & ~x05 & x40 & ~x02 & ~x03))) | (~x04 & ~x05 & ~x02 & ~x03 & x15 & ~x16 & x17 & x40))) | (~x02 & ~x03 & ~x04 & ~x05 & x12 & x40 & (x30 ? (x32 & x33) : ~x31)))) | (~x02 & ~x03 & x12 & ~x13 & (x04 ? (~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : ((~x15 & ((x17 & ((~x19 & (x05 ? (~x16 & (~x18 | (x18 & (x20 ? ~x21 : (x21 & (((x27 | (~x24 & ~x27)) & (~x22 | (x22 & ~x23))) | (x22 & x23 & x27 & (~x24 | (x24 & ~x26))))))))) : (x40 & (x16 ? (~x18 & (~x38 | ~x39)) : (x18 & (x20 ^ x21)))))) | (~x05 & x16 & ~x18 & x19 & x40))) | (~x05 & x16 & x18 & ~x19 & x40))) | (~x05 & x15 & ~x16 & x40 & ((x18 & (~x19 | (~x17 & x19))) | (x17 & ~x18 & x19)))))))) | (~x12 & x13 & ((x01 & ((x16 & (x15 ? (~x17 & ~x18 & ~x19 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))) | (~x02 & (x05 ? ~x03 : x04)))) : (x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))) | (x15 & ~x17 & ~x18 & ((x19 & ((~x02 & ~x03 & ~x04) | (~x16 & ((x02 & (~x03 | (x03 & x04))) | (x03 & ~x04) | (~x02 & x04))))) | (~x02 & ~x03 & ~x04 & ~x05 & ~x19))))) | (x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05)))))))) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x14 & x40 & (x12 ? (x13 ? (~x17 & ((x15 & ~x16 & x18) | (~x18 & ~x19 & ~x15 & x16))) : x15) : x13)));
  assign z08 = ~x08 & ((x09 & (~x10 | (x10 & x11))) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x09 & ~x10 & ~x11 & ~x14 & ~x36 & x40 & ((~x17 & ((x12 & ~x13 & ~x19 & ((~x15 & x16 & x18) | (x15 & ~x16 & ~x18 & ~x37 & ~x38 & ~x39))) | (x15 & ~x16 & ~x12 & x13 & ~x38 & ~x39 & x18 & ~x37))) | (x12 & ~x13 & ~x15 & x16 & x17 & ~x18 & ~x19 & (~x38 | ~x39)))));
  assign z09 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & x40 & ((x13 & (x12 ? ((x14 & x15 & ~x16 & ~x17 & x18) | (~x14 & ~x30)) : (x14 & ~x15))) | (x12 & ~x13 & ~x14 & ~x15 & x16 & ~x19 & (x17 ? (~x18 & (~x38 | ~x39)) : x18)));
  assign z10 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & x40 & ((x12 & ~x13 & ~x14 & ~x15 & x16 & ~x19 & (x17 ? (~x18 & (~x38 | ~x39)) : x18)) | (x13 & (x12 ? ((x14 & x15 & ~x16 & ~x17 & x18) | (~x14 & (~x30 | (x30 & (~x32 | (x32 & ~x33)))))) : (~x15 & (x14 | (~x14 & ~x16))))));
  assign z11 = ~x08 & ((x09 & (~x10 | (x10 & x11))) | (~x01 & ~x02 & ~x03 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x00 & ((~x14 & ((x12 & (x04 ? (~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : ((~x13 & ((~x16 & (x05 ? (~x15 & x17 & x18 & ~x19 & (x20 ? ~x21 : (x21 & (((x27 | (~x24 & ~x27)) & (~x22 | (x22 & ~x23))) | (x22 & x23 & x27 & (~x24 | (x24 & ~x26))))))) : (x15 & ~x18 & x40 & ((x17 & x19) | (~x37 & ~x38 & ~x39 & ~x17 & ~x19))))) | (~x05 & ~x15 & x16 & x19 & x40 & x17 & ~x18))) | (~x05 & x13 & x40 & (~x30 | (x30 & (~x32 | (x32 & (~x33 | (x33 & x35)))))))))) | (~x04 & ~x12 & x13 & ((~x05 & x40 & ((x15 & ~x17 & (~x18 | (~x16 & x18 & ~x37 & ~x38 & ~x39))) | (x17 & x18 & x19 & ~x15 & x16))) | (x17 & ~x18 & ~x19 & x05 & ~x15 & x16))))) | (~x04 & ~x05 & x12 & x13 & x14 & x15 & ~x16 & ~x17 & x18 & x40))) | (~x05 & x12 & ~x13 & x00 & ~x04 & x17 & ~x18 & ~x19 & ~x14 & ~x15 & ~x16))));
  assign z12 = ~x01 & ~x02 & ~x03 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x05 & x12 & ~x13 & x00 & ~x04 & x17 & ~x18 & ~x19 & ~x14 & ~x15 & ~x16) | (~x00 & ((~x04 & ~x05 & x12 & x13 & x14 & x15 & ~x16 & ~x17 & x18 & x40) | (~x14 & ((~x04 & ~x12 & x13 & ((~x05 & x40 & ((x15 & ~x17 & (~x18 | (~x16 & x18 & ~x37 & ~x38 & ~x39))) | (x17 & x18 & x19 & ~x15 & x16))) | (x17 & ~x18 & ~x19 & x05 & ~x15 & x16))) | (x12 & (x04 ? (~x05 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : ((~x13 & ((~x16 & (x05 ? (~x15 & x17 & x18 & ~x19 & (x20 ? ~x21 : (x21 & (((x27 | (~x24 & ~x27)) & (~x22 | (x22 & ~x23))) | (x22 & x23 & x27 & (~x24 | (x24 & ~x26))))))) : (x15 & ~x18 & x40 & ((x17 & x19) | (~x37 & ~x38 & ~x39 & ~x17 & ~x19))))) | (~x05 & ~x15 & x16 & x19 & x40 & x17 & ~x18))) | (~x05 & x13 & x40 & (~x30 | (x30 & (~x32 | (x32 & (~x33 | (x33 & x35)))))))))))))));
  assign z13 = ~x08 & ((x09 & (~x10 | (x10 & x11))) | (~x01 & ~x02 & ~x03 & ~x09 & ~x10 & ~x11 & ~x14 & ~x36 & ((~x00 & (x04 ? (x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : (x05 ? (~x15 & x17 & ~x19 & ((x12 & ~x13 & ~x16 & x18 & (x20 ? ~x21 : (x21 & (((x27 | (~x24 & ~x27)) & (~x22 | (x22 & ~x23))) | (x22 & x23 & x27 & (~x24 | (x24 & ~x26))))))) | (~x12 & x13 & x16 & ~x18))) : (x40 & ((x13 & (x12 ? (~x30 | (x30 & (~x32 | (x32 & (~x33 | (x33 & x35)))))) : ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18)))) | (x12 & ~x13 & ((x17 & ~x18 & ((x19 & (x15 ^ x16)) | (~x15 & x16 & ~x19 & (~x38 | ~x39)))) | (~x15 & x16 & ~x17 & x18 & ~x19)))))))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & ~x05 & x12 & ~x13 & x00 & ~x04))));
  assign z14 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x02 & (x00 ? (~x01 & ~x04 & ~x05 & ~x14 & ((~x12 & x13 & ((x16 & ((x03 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x03 & x15 & ~x17 & ~x18 & x19))) | (~x17 & ~x18 & ~x19 & ~x03 & x15 & ~x16))) | (~x16 & x17 & ~x18 & ~x19 & ~x13 & ~x15 & ~x03 & x12))) : ((~x14 & ((~x03 & ((~x18 & ((~x12 & x13 & ((~x17 & ((x01 & x15 & ((x04 & ~x05 & x16 & x19) | (~x16 & ~x19 & ~x04 & x05))) | (~x01 & ~x04 & ~x05 & ~x15 & x16 & ~x19 & x40))) | (~x01 & ~x04 & ~x15 & x16 & x17 & (x05 ? ~x19 : (x19 & x40))))) | (~x01 & ~x04 & ~x05 & x12 & ~x13 & x40 & ((~x16 & (x15 ? (x19 | (x17 & ~x19)) : (x17 & x19 & (~x37 | x38 | ~x39)))) | (~x15 & x16 & x17 & (x19 | (~x19 & (~x38 | ~x39)))))))) | (~x01 & ((x12 & ((~x13 & ((x18 & ((~x16 & ((~x04 & ~x19 & ((x05 & ~x15 & x17 & x20 & x21) | (~x05 & x15 & x40))) | (x04 & x05 & x15 & ~x17 & x19))) | (~x04 & ~x05 & ~x15 & x40 & ((x17 & x19) | (x16 & (~x17 ^ ~x19)))))) | (~x04 & ~x05 & ~x15 & ~x17 & x40 & (~x16 | (x16 & ~x19))))) | (~x04 & ~x05 & x13 & x40 & (~x15 | (x15 & ~x16))))) | (~x04 & ~x05 & ~x12 & x13 & x40 & ((~x15 & (~x16 | (x16 & (x19 ? ~x17 : x18)))) | (x17 & x18 & x19 & x15 & ~x16))))))) | (~x01 & x03 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x19 & ((x18 & ((~x20 & x21 & ((~x05 & (((x22 ? (x23 & ~x24) : x24) & (~x04 ^ x27)) | (~x04 & x22 & x24 & ~x27 & (~x23 | (x23 & ~x25))))) | (~x04 & x05 & (x22 ? ((x24 & (x27 | (x23 & x25 & ~x27))) | (~x23 & ~x24 & ~x27)) : (~x24 & ~x27))))) | (~x04 & x05 & x20 & ~x21 & ~x27))) | (~x04 & ~x05 & ~x18))))) | (~x01 & ~x03 & ~x04 & ~x05 & x14 & x40 & (x12 ? (~x13 | (x13 & ((~x16 & ((~x17 & ((x18 & ~x19) | (x15 & (~x18 | (x18 & x19))))) | (~x15 & (x18 ? x17 : x19)))) | (~x17 & ~x19 & (x15 ? x16 : ~x18))))) : (x13 | (~x16 & ~x17 & x18 & ~x13 & ~x15))))))) | (~x00 & ~x01 & x02 & ~x03 & ~x04 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x05 ? (x20 & ~x21) : (~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))));
  assign z15 = (~x08 & (x09 ? (~x10 | (x10 & x11)) : (x10 | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x10 & ~x11 & ~x36 & x40 & ((x15 & ((~x14 & (x05 ? (x12 & ~x13 & (x17 ? ((x18 & x19) | (x16 & (~x18 | (x18 & ~x19)))) : x16)) : ((~x12 & x13 & ((x16 & (x18 | (x17 & ~x18))) | (~x16 & ~x17 & x18 & ~x38 & ~x39))) | (~x16 & ~x17 & x12 & ~x13 & ~x18 & ~x19 & ~x38 & ~x39)))) | (x05 & x14 & ((x17 & (x12 ? (x13 & (~x16 | (x16 & x18 & ~x19))) : (~x13 & x16))) | (~x12 & ~x13 & ~x16))))) | (~x13 & ((~x12 & (x05 ? (x14 & (x17 ? ~x15 : x16)) : ~x14)) | (~x14 & ~x15 & ~x16 & ~x05 & x12 & x17 & ~x18 & x19 & x37 & ~x38))) | (x05 & x12 & x13 & x14 & x16 & ((~x15 & (x19 ? ~x17 : x18)) | (x17 & (~x18 | (x18 & x19)))))))))) | (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36);
  assign z16 = ~x08 & (x09 ? x10 : (~x10 & ~x11 & (x36 | (~x36 & (x00 ? (~x01 & ~x02 & ~x03 & ~x12 & x13 & ~x14 & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18 & ((x16 & ~x19) | (~x16 & x19 & ~x04 & ~x05))))) : ((~x14 & ((~x12 & x13 & ((x01 & ((x16 & (x15 ? (~x17 & ~x18 & ~x19 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))) | (~x02 & (x05 ? ~x03 : x04)))) : (x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))) | (x15 & ~x17 & ~x18 & ((x19 & ((~x02 & ~x03 & ~x04) | (~x16 & ((x02 & (~x03 | (x03 & x04))) | (x03 & ~x04) | (~x02 & x04))))) | (~x02 & ~x03 & ~x04 & ~x05 & ~x19))))) | (x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))))) | (~x01 & ((~x02 & ((~x16 & (x12 ? (~x13 & ((~x19 & ((~x15 & x17 & ((x18 & (x03 ? ((x27 & ((((x20 & ~x21) | (~x20 & x21 & x22 & ~x23 & ~x24)) & (x05 | (x04 & ~x05))) | (~x20 & x21 & (x04 ? (~x22 & ~x24) : (~x22 | (x22 & ((x23 & ~x24) | (~x05 & (~x23 | (x23 & x24)))))))))) | (~x04 & ~x05 & (x20 ? ~x21 : (x21 & ~x27 & (x22 ? (x23 ? (x24 & x25) : ~x24) : ~x24))))) : (((x20 ^ x21) & (x05 | (x04 & ~x05))) | (~x04 & ~x05 & x40 & (x20 | (~x20 & x21)))))) | (~x03 & ~x18 & (x05 | (~x05 & (x04 | (~x04 & x40))))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18 & x40 & (x38 | x39 | (~x37 & ~x38 & ~x39))))) | (~x03 & x19 & ((x15 & x18 & (x04 ? (~x05 & ~x17) : (x05 ? ~x17 : x40))) | (~x04 & ~x05 & ~x15 & x17 & ~x18 & x39 & x40))))) : (x13 & x15 & ((~x03 & ((x17 & (((x05 | (x04 & ~x05)) & (~x19 | (~x18 & x19))) | (~x04 & ~x05 & ~x19 & x40))) | (~x04 & ~x05 & x40 & ((~x18 & x19) | (~x17 & x18 & (x38 | x39 | (~x37 & ~x38 & ~x39))))))) | (x03 & ~x04 & ~x05 & x17 & ~x18))))) | (~x12 & x13 & (((x05 ? ~x03 : x04) & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18))) | (~x03 & ~x04 & ~x05 & x40 & ((x17 & x18 & x19 & ~x15 & x16) | (~x18 & ((x15 & ~x17 & (~x19 | (x16 & x19))) | (x17 & ~x19 & ~x15 & x16))))))) | (~x03 & ~x04 & ~x05 & x12 & ~x13 & x16 & x40 & (x15 | (~x15 & x17 & ~x18 & ~x19 & (x38 | x39)))))) | (x02 & ((~x03 & ((~x12 & x13 & x15 & ~x17 & ~x18) | (~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x20 & ~x21 & x27))) | (x03 & x04 & ~x05 & ~x12 & x13 & x15 & ~x17 & ~x18))) | (x03 & ~x12 & x13 & (~x04 | (x04 & x05)) & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18))))))) | (~x01 & ~x02 & ~x03 & ~x04 & ~x05 & (~x40 | (x14 & x40 & ((x16 & ((x17 & (x12 ? (x13 & (~x18 | (x18 & (x19 | (x15 & ~x19))))) : (~x13 & (~x18 | (x15 & x18))))) | (x12 & x13 & ~x15 & (x19 ? ~x17 : x18)) | (~x12 & ~x13 & ~x17))) | (~x16 & ((~x12 & ~x13 & (x15 | (~x15 & ~x18))) | (x12 & x13 & x15 & x17))) | (~x12 & ~x13 & ~x15 & x17 & x18)))))))))));
  assign z17 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & x40 & ((~x15 & ((x12 & ((x13 & x14 & ~x16 & (x17 ? (~x18 & ~x19) : (x18 & x19))) | (~x17 & ~x18 & x19 & ~x13 & ~x14 & x16))) | (~x12 & ~x13 & x14 & ~x16 & ~x17 & ~x18))) | (x12 & x13 & x15 & x16 & (~x14 | (x14 & ~x17 & x19))));
  assign z18 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & (x09 ? (~x10 | (x10 & x11)) : (x10 | (~x00 & ~x01 & ~x02 & ~x04 & ~x05 & ~x10 & ~x11 & ~x16 & ~x36 & ((x13 & ((~x12 & ~x14 & x15 & ((x03 & x17 & (~x19 | (~x18 & x19))) | (~x03 & ~x17 & x18 & x37 & ~x38 & ~x39 & x40))) | (~x03 & x12 & x14 & ~x15 & x40 & (x17 ? (~x18 & ~x19) : (x18 & x19))))) | (~x03 & ~x13 & ~x18 & x40 & ((x12 & ~x14 & x37 & ~x38 & ((~x15 & x17 & x19) | (x15 & ~x17 & ~x19 & ~x39))) | (~x12 & x14 & ~x15 & ~x17))))))));
  assign z19 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & (x10 ? x11 : (x09 | (~x00 & ~x01 & ~x02 & ~x04 & ~x09 & ~x11 & ~x36 & ((~x05 & ((~x14 & ((~x12 & ((x15 & ((x13 & ((~x16 & ((x03 & x17 & (~x19 | (~x18 & x19))) | (~x03 & ~x17 & x18 & ~x38 & ~x39 & x40))) | (~x03 & x16 & x18 & x40 & (~x17 | (x17 & ~x19))))) | (~x03 & x40 & ((~x13 & (~x16 | (x16 & ~x17))) | (x16 & x17 & (~x18 | (x18 & x19))))))) | (~x03 & ~x13 & x40 & ((x17 & ((~x15 & ~x18) | (x16 & x18 & ~x19))) | (~x15 & (x16 ? (x19 ? x18 : ~x17) : x18)))))) | (~x03 & x40 & ((x12 & (x13 ? (x15 & x16) : (~x16 & ~x18 & ~x38 & ((x15 & ~x17 & ~x19 & ~x39) | (~x15 & x17 & x19 & x37))))) | (~x17 & ~x18 & x19 & ~x13 & ~x15 & x16))))) | (~x03 & x40 & ((~x15 & ~x16 & ((x12 & x13 & x14 & (x17 ? (~x18 & ~x19) : (x18 & x19))) | (~x17 & ~x18 & ~x12 & ~x13))) | (x12 & x13 & x14 & ~x17 & x19 & x15 & x16))))) | (~x03 & x05 & x40 & ((x14 & ((x15 & ((x17 & (x12 ? (x13 & (~x16 | (x16 & x18 & ~x19))) : (~x13 & x16))) | (~x12 & ~x13 & ~x16))) | (~x12 & ~x13 & (x17 ? ~x15 : x16)) | (x12 & x13 & x16 & ((~x15 & (x19 ? ~x17 : x18)) | (x17 & (~x18 | (x18 & x19))))))) | (x12 & ~x13 & ~x14 & x15 & (x17 ? ((x18 & x19) | (x16 & (~x18 | (x18 & ~x19)))) : x16)))))))));
  assign z20 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & (x00 ? (~x01 & ~x02 & ~x12 & x13 & ~x14 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))) : ((~x01 & ((~x04 & (x03 ? (~x14 & ((~x12 & x13 & x15 & ~x17 & ~x18) | (~x15 & x17 & x18 & ((~x02 & x12 & ~x13 & ~x16 & ~x19 & ((~x20 & x21 & (x27 ? ((x05 & (x22 ? (x23 & (~x24 | (x24 & ~x26))) : x24)) | (x22 & x23 & x24 & x26)) : (x05 ? ((~x22 & ~x24) | (x24 & x25 & x22 & x23)) : (x22 ? x23 : x24)))) | (~x21 & ~x27 & x05 & x20))) | (x16 & x19 & ~x12 & x13))))) : ((x12 & ((~x14 & ((~x13 & ((x17 & ((~x19 & ((~x15 & (x02 ? (~x16 & x18 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x22 & ~x24))) : (~x05 & x16 & ~x18 & x40 & (~x38 | ~x39)))) | (~x02 & ~x05 & x15 & x40 & (~x18 | (x16 & x18))))) | (~x02 & ~x05 & x19 & x40 & (x18 | (x15 & x16 & ~x18))))) | (~x02 & ~x05 & x40 & (x15 ? (~x17 & ((x16 & (~x18 | (x18 & x19))) | (~x16 & x19) | (x18 & ~x19))) : (x16 ? (~x17 & x18) : (~x18 & ~x19)))))) | (~x02 & ~x05 & x13 & ~x15 & x40 & ((x20 & x21 & x29) | (~x29 & ~x31))))) | (~x02 & ~x05 & x14 & x40 & (x13 ? ((x15 & ((~x16 & (~x18 | (x17 & x18))) | (x18 & ~x19 & x16 & x17))) | (~x18 & ((x16 & x17) | (~x15 & ~x17 & ~x19))) | (~x15 & ((x16 & ~x17 & (x19 | (x18 & ~x19))) | (x17 & (x19 ? ~x16 : x18)))) | (x18 & x19 & x16 & x17)) : ~x15)))) | (~x02 & ~x12 & ((~x05 & x40 & ((x14 & (x13 | (~x13 & ((~x16 & (x15 | (~x15 & x18 & x19))) | (x16 & ~x17) | (x17 & (((~x18 | (x18 & ~x19)) & (~x15 | (x15 & x16))) | (x16 & x18 & x19))))))) | (x13 & ~x14 & ((x17 & ((~x15 & x16 & ~x18) | (x18 & x19 & x15 & ~x16))) | (~x17 & ~x18 & ((x16 & ~x19) | (x15 & (~x16 | (x16 & x19))))) | (~x15 & (~x16 | (x16 & x18 & x19))))))) | (~x14 & ~x15 & x05 & x13 & ~x18 & ~x19 & x16 & x17)))))) | (~x14 & ((~x12 & x13 & (x15 ? (~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (~x02 & (x05 ? ~x03 : x04)) | (x03 & x04 & x05))) : (x16 & x17 & x18 & x19 & ((~x02 & (x05 ? ~x03 : x04)) | (x03 & x04 & x05))))) | (~x02 & x03 & x04 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & ~x20 & x21 & x27 & (x05 ? (~x22 & ~x24) : (x22 ? (x23 & ~x24) : x24))))))) | (~x12 & x13 & ~x14 & ((x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))) | (x01 & (x15 ? (~x17 & ~x18 & ((x04 & ((((~x16 & x19) | (x05 & x16 & ~x19)) & (~x02 | (x02 & x03))) | (~x05 & x16 & (x03 ? ~x19 : ~x02)))) | (~x02 & ~x03 & ~x04) | ((~x16 ^ ~x19) & (x03 ? ~x04 : x02)))) : (x16 & x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05)))))))))));
  assign z21 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x14 & x15 & ~x16 & ~x36 & x40 & ((~x12 & x13 & x17 & (~x19 | (~x18 & x19))) | (x12 & ~x13 & ~x17 & x18));
  assign z22 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & (x10 | (~x10 & (x09 | (~x09 & ~x11 & (x36 | (~x01 & ~x36 & ((~x00 & ((~x02 & ((~x04 & ((~x05 & ((~x14 & ((~x13 & ((~x19 & ((x12 & (x03 ? (~x15 & ~x16 & x17 & (~x18 | (x18 & (x20 ? ~x21 : (x21 & (x22 ? (x24 ? (~x23 | (x23 & ~x26 & x27)) : x27) : (x27 | (~x24 & ~x27)))))))) : (x40 & ((~x18 & (((x38 | x39) & (x15 ? (~x16 & ~x17) : (x16 & x17))) | (x15 & ~x16 & ~x17 & ~x38 & ~x39))) | (~x16 & x18 & (x15 | (~x15 & x17 & (x20 | (~x20 & x21))))))))) | (~x03 & x40 & ((~x12 & ((x15 & ((~x17 & x18) | (~x16 & x17 & ~x18))) | (x16 & (x17 ? ~x18 : ~x15)) | (~x16 & x17 & x18))) | (~x15 & x16 & x17 & x18))))) | (~x03 & x40 & (x15 ? ((~x12 & (x17 ? (x18 & x19) : ~x18)) | (~x16 & x19 & (x17 ^ x18))) : ((~x12 & ((x18 & x19) | (~x16 & x17 & ~x18))) | (~x18 & ((x12 & (x16 ? ~x17 : x19)) | (x16 & x17 & x19))) | (~x17 & x18 & x12 & ~x16)))))) | (~x12 & ((x15 & ((x13 & ((~x16 & (x03 ? (x17 & (~x19 | (~x18 & x19))) : (~x17 & x18 & x40 & (x38 | x39 | (~x38 & ~x39))))) | (~x03 & x16 & x40 & (x17 ? (~x18 ^ x19) : (x18 & ~x19))))) | (~x03 & x16 & x40 & (x17 ? (x18 ^ x19) : (x18 & x19))))) | (~x03 & ~x15 & x16 & x40 & ((~x17 & ~x18 & x19) | (x13 & x18 & ~x19))))) | (~x03 & x12 & x13 & x40 & (x15 | (~x15 & ~x29))))) | (~x03 & (~x40 | (x40 & ((~x16 & ((~x17 & ((~x15 & ((~x12 & ~x13 & (~x19 | (~x18 & x19))) | (x12 & x13 & x14 & ~x18 & x19))) | (x12 & x13 & x14 & (x18 | (x15 & ~x18))))) | (x12 & x13 & x14 & ~x18 & ~x19 & ~x15 & x17))) | (x14 & x15 & (x12 ? (~x13 | (x13 & x16 & ~x17)) : x13)))))))) | (x05 & ((x12 & ((x17 & ((x18 & ((~x13 & ~x14 & ((~x19 & ((~x15 & ~x16 & (x03 ? (~x20 & x21 & x27 & (x22 ? ~x23 : ~x24)) : x20)) | (x16 & x40 & ~x03 & x15))) | (x19 & x40 & ~x03 & x15))) | (~x03 & x13 & x14 & x16 & x40 & (x19 | (x15 & ~x19))))) | (~x03 & x40 & ((x13 & x14 & (x16 ? ~x18 : x15)) | (x15 & x16 & ~x18 & ~x13 & ~x14))))) | (~x03 & x16 & x40 & ((x13 & x14 & ~x15 & (x19 ? ~x17 : x18)) | (x15 & ~x17 & ~x13 & ~x14))))) | (~x03 & ~x12 & ~x13 & x14 & x40 & ((~x15 & x17) | (x16 & ~x17) | (x15 & (~x16 | (x16 & x17))))))) | (x03 & x12 & ~x13 & ~x16 & x17 & ~x14 & ~x15 & x18 & ~x19 & ~x20 & x21 & ~x24 & ~x27 & x22 & ~x23))) | (~x14 & ~x16 & (((x05 | (x04 & ~x05)) & ((~x03 & ((x17 & ((~x19 & (x12 ? (~x13 & ~x15 & (~x18 | (x18 & ~x20 & x21))) : (x13 & x15))) | (~x12 & x13 & x15 & ~x18 & x19))) | (~x17 & x18 & x19 & x12 & ~x13 & x15))) | (x03 & x12 & ~x13 & ~x15 & x17 & x18 & ~x19 & x20 & ~x21 & x27))) | (x04 & x12 & ~x13 & ~x15 & x17 & x18 & ~x19 & (x03 ? (~x20 & x21 & ~x24 & x27 & (x22 ? ~x23 : ~x05)) : (x20 & ~x21))))))) | (~x04 & ~x05 & x02 & ~x03 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & ~x20 & x21 & x22 & ~x23 & ~x24 & x27))) | (~x04 & ~x05 & x12 & x00 & ~x02 & ~x03 & ~x16 & x17 & ~x18 & ~x19 & ~x13 & ~x14 & ~x15)))))))));
  assign z23 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & x40 & ((x13 & ((x14 & x15 & (~x12 | (~x17 & ~x18 & x12 & ~x16))) | (x12 & ~x14 & ~x15 & (~x29 | (x29 & (~x20 | (x20 & ~x21))))))) | (x12 & ~x13 & ~x14 & x15 & ~x16 & ~x17 & x18));
  assign z24 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & (x10 | (~x10 & (x09 | (~x09 & ~x11 & (x36 | (~x36 & (x00 ? (~x01 & ~x02 & ~x14 & ((~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x12 & x13 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))))) : ((~x01 & ((~x02 & ((~x14 & ((~x04 & ((~x13 & ((x17 & ((~x19 & ((~x15 & ((x12 & ((~x05 & (x03 ? (~x16 & (~x18 | (x18 & ~x20 & x21 & x22 & (x24 ? ~x23 : x27)))) : (x40 & (x16 ? (~x18 & (x38 | x39)) : (x18 & (x20 | (~x20 & x21))))))) | (~x16 & x18 & ((x20 & (x03 ? ~x21 : x05)) | (x03 & ~x20 & x21 & (x22 ? ((~x23 & ~x24 & ~x27) | (x27 & ((x05 & (~x23 | (x23 & ~x24))) | (x23 & x24 & ~x26)))) : (x27 | (~x24 & ~x27)))))))) | (~x03 & ~x05 & x18 & x40 & (x16 | (~x12 & ~x16))))) | (~x03 & x40 & ((~x05 & ((x15 & ~x16 & x18) | (~x12 & ~x18 & (x16 | (x15 & ~x16))))) | (x05 & x12 & x15 & x16 & x18))))) | (~x03 & x40 & ((x15 & (x05 ? (x12 & (x18 ? x19 : x16)) : (~x16 & x19 & (~x18 | (~x12 & x18))))) | (~x05 & ((~x12 & ((~x15 & ~x16 & ~x18) | (x16 & x18 & x19))) | (~x18 & x19 & ~x15 & x16))))))) | (~x03 & x40 & ((~x05 & ((~x17 & (x15 ? ((~x19 & (x12 ? (~x16 & ~x18 & (x38 | x39 | (~x38 & ~x39))) : (x18 | (x16 & ~x18)))) | (~x12 & ~x16 & x19)) : ((x16 & (~x18 | (~x12 & x18))) | (x12 & ~x16 & x18)))) | (~x15 & ~x16 & x19 & (x12 ^ x18)))) | (x05 & x12 & x15 & x16 & ~x17))))) | (~x05 & ((~x12 & ((x15 & ((x13 & ((~x03 & x16 & x40 & (x17 ? (~x18 ^ x19) : (x18 & ~x19))) | (~x16 & ((~x03 & ~x17 & x18 & x40 & (x38 | x39 | (~x38 & ~x39))) | (x17 & (x03 ? (~x19 | (~x18 & x19)) : x40)))))) | (~x03 & x40 & ((x16 & (x17 ? (x18 ^ x19) : x19)) | (~x18 & ~x19 & ~x16 & ~x17))))) | (~x03 & x13 & ~x15 & x16 & x40 & (~x18 | (x18 & ~x19))))) | (~x03 & x12 & x13 & x40 & (x15 | (~x15 & x20 & x21 & ~x22 & x23 & x29))))))) | (~x16 & ((x17 & (x03 ? (x04 & x12 & ~x13 & ~x15 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : (((x05 | (x04 & ~x05)) & ((~x12 & x13 & x15 & ~x18 & x19) | (x12 & ~x13 & ~x15 & ~x19 & (~x18 | (x18 & ~x20 & x21))))) | (~x19 & ((x04 & ((x13 & x15 & ~x05 & ~x12) | (x12 & ~x13 & ~x15 & x18 & x20 & ~x21))) | (x05 & ~x12 & x13 & x15 & x18)))))) | (x15 & ((~x17 & ((~x03 & x12 & ~x13 & x18 & x19 & (x05 | (x04 & ~x05))) | (x04 & ~x05 & ~x12 & x13 & ~x18 & ~x19))) | (x13 & ~x18 & ~x19 & ~x03 & x05 & ~x12))))) | (~x12 & x13 & x16 & ((x04 & ((x18 & x19 & ~x15 & x17) | (x15 & ~x17 & ~x18 & (~x19 | (~x05 & x19))))) | (~x17 & ~x18 & x19 & ~x03 & x05 & x15))))) | (~x03 & ~x04 & (x40 ? ((x14 & ((x12 & ((x13 & (x05 ? ((x17 & ((x16 & (~x18 | (x18 & x19))) | (x15 & (~x16 | (x16 & x18 & ~x19))))) | (~x15 & x16 & (x19 ? ~x17 : x18))) : ((~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x17 & ((x15 & (x16 | (~x16 & ~x18))) | (~x16 & (x18 | (~x15 & ~x18 & x19)))))))) | (~x05 & ~x13 & x15))) | (x05 & ~x12 & ~x13 & ((~x15 & x17) | (x16 & ~x17) | (x15 & (~x16 | (x16 & x17))))))) | (~x05 & ~x12 & ~x13 & ~x15 & ~x16 & ~x17 & (~x19 | (~x18 & x19)))) : ~x05)))) | (~x14 & ((~x12 & x13 & ((x15 & ~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05 & (~x16 ^ x19)))))) | (x18 & x19 & x16 & x17 & x03 & ~x04 & ~x15))) | (x02 & ~x03 & ~x04 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))))))) | (~x12 & x13 & ~x14 & ((x16 & ((x01 & (x15 ? (~x17 & ~x18 & ~x19 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (~x02 & (x05 ? ~x03 : x04)) | (x03 & (~x04 | (~x02 & x04 & x05))))) : (x17 & x18 & x19 & (~x02 | (x02 & x03 & ~x04))))) | (x02 & ((x03 & x04 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))) | (x17 & x18 & x19 & ~x03 & ~x15))))) | (x15 & ~x17 & ~x18 & ((x01 & ((~x02 & ~x03 & ~x04 & ~x05 & ~x19) | (x19 & ((~x02 & ~x03 & ~x04) | (~x16 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & ~x04))))))) | (x04 & ~x16 & x19 & (~x02 | (x02 & x03 & x05))))))))))))))));
  assign z25 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & (x00 ? (~x01 & ~x02 & ~x12 & x13 & ~x14 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))) : ((x13 & ((~x18 & ((~x17 & ((~x02 & ((~x01 & ((~x12 & ~x14 & ((x15 & ((((x04 & ~x05) | (~x03 & (x05 | (~x04 & ~x05 & x40)))) & (~x16 ^ x19)) | (x04 & x16 & ~x19))) | (~x03 & ~x04 & ~x05 & ~x15 & x16 & ~x19 & x40))) | (~x03 & ~x04 & ~x05 & x12 & x14 & ~x16 & x40 & (x15 | (~x15 & x19))))) | (~x12 & ~x14 & x15 & ((x01 & ((~x19 & ((~x03 & (x05 ? x16 : ~x04)) | (x04 & x16 & (~x05 | (x03 & x05))))) | (~x03 & ~x04 & x19))) | (x04 & ~x16 & x19))))) | (~x12 & ~x14 & x15 & (((~x16 ^ ~x19) & ((x02 & ((x03 & x04 & x05) | (x01 & (~x03 | (x03 & x04 & ~x05))))) | (x01 & x03 & ~x04))) | (~x01 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05 & (~x16 ^ x19)))))))))) | (~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x12 & ~x14 & ~x15 & x16 & x17 & x40))) | (~x14 & ((~x15 & ((~x12 & x16 & x17 & x18 & x19 & ((x01 & (~x02 | (x02 & x03 & ~x04))) | (x02 & (~x03 | (x03 & x04))) | (~x01 & (x04 ? ~x02 : x03)))) | (~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x12 & x40 & (~x29 | (x29 & (~x20 | (x20 & (~x21 | (x21 & ~x22 & x23))))))))) | (~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x12 & x18 & x19 & x40 & x15 & ~x16 & x17))))) | (~x01 & ~x04 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & ((x27 & (x02 ? (~x03 & ((x05 & x20 & ~x21) | (~x05 & ~x20 & x21 & ~x22 & ~x24))) : (x03 & x05 & ~x20 & x21 & (x22 ? (x23 & (~x24 | (x24 & ~x26))) : x24)))) | (~x02 & x03 & x05 & ~x27 & ((x20 & ~x21) | (~x20 & x21 & ~x22 & ~x24)))))));
  assign z26 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & (x00 ? (~x01 & ~x02 & ~x03 & ~x12 & x13 & ~x14 & ((x16 & (x04 ? (~x05 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) : ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15)))) | (~x04 & ~x05 & x15 & ~x17 & ~x18))) : ((~x01 & ((~x04 & (x12 ? ((~x14 & ((~x02 & (x03 ? (x05 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & (x20 ? (~x21 & ~x27) : (x21 & (x22 ? (x23 & (x27 | (x24 & x25 & ~x27))) : (x24 ^ ~x27))))) : (~x05 & x40 & ((~x15 & (x13 ? (x20 & x21 & x29 & (x23 | (x22 & ~x23))) : ((~x16 & x17 & ~x18 & ~x19) | (x16 & (x17 ? (~x18 & ~x19 & (~x38 | ~x39)) : x18))))) | (~x13 & x15 & ((x18 & ((x16 & (~x17 ^ ~x19)) | (x17 & x19) | (~x17 & ~x19))) | (x16 & ~x18) | (~x16 & ~x17 & x19))))))) | (x17 & x18 & ~x19 & x20 & ~x21 & x27 & ~x13 & ~x15 & ~x16 & x02 & ~x03 & ~x05))) | (~x02 & ~x03 & ~x05 & x14 & x40 & (x13 ? ((x17 & ((x15 & (~x16 | (x16 & x18 & ~x19))) | (x16 & (~x18 | (x18 & x19))) | (~x15 & x18 & ~x19))) | (~x15 & (x16 ? (~x17 & (x19 | (x18 & ~x19))) : (~x18 & x19)))) : ~x15))) : ((x13 & ((~x14 & ((x03 & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18))) | (~x02 & ~x03 & ~x05 & x40 & ((x17 & ((~x15 & x16 & ~x18) | (x18 & x19 & x15 & ~x16))) | (~x17 & ~x18 & ((x16 & ~x19) | (x15 & (~x16 | (x16 & x19))))) | (~x15 & (~x16 | (x16 & x18 & x19))))))) | (~x02 & ~x03 & ~x05 & x14 & ~x15 & x40))) | (~x02 & ~x03 & ~x05 & ~x13 & x14 & x40 & ((~x16 & (x15 | (~x15 & x18 & x19))) | (x16 & ~x17) | (x17 & (((~x18 | (x18 & ~x19)) & (~x15 | (x15 & x16))) | (x16 & x18 & x19)))))))) | (~x14 & ((~x12 & x13 & (x15 ? (~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (~x02 & (x05 ? ~x03 : x04)) | (x03 & x04 & x05))) : (x16 & x17 & x18 & x19 & ((~x02 & (x05 ? ~x03 : x04)) | (x03 & x04 & x05))))) | (x04 & x05 & ~x02 & x03 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & ~x20 & ~x24 & x27 & x21 & ~x22))))) | (~x12 & x13 & ~x14 & ((x01 & ((x16 & (x15 ? (~x17 & ~x18 & ~x19 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))) | (~x02 & (x05 ? ~x03 : x04)))) : (x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))) | (x15 & ~x17 & ~x18 & ((x19 & ((~x02 & ~x03 & ~x04) | (~x16 & ((x02 & (~x03 | (x03 & x04))) | (x03 & ~x04) | (~x02 & x04))))) | (~x02 & ~x03 & ~x04 & ~x05 & ~x19))))) | (x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05)))))));
  assign z27 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & ((x10 & (~x09 | (x09 & ~x11))) | (~x09 & ~x10 & ~x11 & (x36 | (~x36 & (x00 ? (~x01 & ~x02 & ~x14 & ((~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x12 & x13 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))))) : ((~x12 & x13 & ~x14 & ((x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))) | (x01 & (x15 ? (~x17 & ~x18 & ((x04 & ((((~x16 & x19) | (x05 & x16 & ~x19)) & (~x02 | (x02 & x03))) | (~x05 & x16 & (x03 ? ~x19 : ~x02)))) | (~x02 & ~x03 & ~x04) | ((~x16 ^ ~x19) & (x03 ? ~x04 : x02)))) : (x16 & x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))))) | (~x01 & ((~x02 & ((~x14 & ((~x13 & ((~x16 & ((x12 & ((~x19 & ((~x15 & ((x17 & (x18 ? (x20 ? ((~x21 & (x03 ? (~x04 | (x04 & x27)) : x04)) | (~x03 & ~x04 & (x05 | (~x05 & x40)))) : (x21 & (x03 ? (x05 ? ((~x24 & (~x22 | (x22 & ~x23)) & (~x04 ^ x27)) | (~x04 & (x27 | (x22 & x23 & x24 & x25 & ~x27)))) : (~x04 | (x04 & x27 & (~x22 | (x22 & ~x24))))) : (x05 | (~x05 & (x04 | (~x04 & x40))))))) : (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05))))) | (~x03 & ~x04 & ~x05 & ~x18 & x40))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18 & x40 & (x38 | x39 | (x37 & ~x38 & ~x39))))) | (~x03 & ((~x05 & ((x19 & ((~x04 & ~x18 & x40 & (x15 | (~x15 & x17))) | (~x17 & x18 & x04 & x15))) | (~x17 & x18 & x40 & ~x04 & ~x15))) | (~x17 & x18 & x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x40 & ((~x12 & ((x17 & (x15 ? x19 : ~x18)) | (~x15 & (x19 ? x18 : ~x17)))) | (~x17 & x19 & (x15 ^ ~x18)) | (x15 & ~x19 & (x18 | (x17 & ~x18))))))) | (~x03 & ~x04 & x40 & ((x16 & ((~x05 & ((~x15 & ((x12 & ~x19 & (x18 | (x17 & ~x18))) | (x17 & ~x18 & x19) | (~x17 & (~x18 | (x18 & x19))))) | (~x12 & (x17 ? (~x18 ^ x19) : (x18 ? ~x19 : x15))))) | (x12 & x15 & (~x17 | (x17 & (~x18 | (x18 & ~x19))))))) | (x17 & x18 & ((~x05 & ~x15 & (~x12 ^ x19)) | (x12 & x15 & x19))))))) | (~x12 & ((x13 & ((x15 & ((~x16 & ((x17 & (((~x19 | (~x18 & x19)) & (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05)))) | (~x05 & x40 & ~x03 & ~x04))) | (~x03 & ~x04 & ~x05 & ~x17 & x18 & x40 & (x38 | x39 | (x37 & ~x38 & ~x39))))) | (~x17 & ~x18 & (x05 ? ~x03 : x04)))) | (~x03 & ((~x15 & ((~x04 & ((x17 & ~x18 & ~x19 & x05 & x16) | (~x05 & ~x16 & x40))) | (x17 & x18 & x19 & x05 & x16))) | (~x04 & ~x05 & x16 & x40))) | (x18 & x19 & x16 & x17 & x04 & ~x05 & ~x15))) | (~x03 & ~x04 & ~x05 & x15 & ~x18 & x40 & ~x16 & ~x17))) | (~x03 & ~x04 & ~x05 & x12 & x13 & x40))) | (~x03 & ~x04 & (x40 ? ((x14 & ((x16 & (x12 ? (x13 & ((x19 & (x05 ? (x17 ? x18 : ~x15) : (x18 & (~x15 | (x15 & x17))))) | (~x05 & ~x17 & (x15 | (~x15 & ~x18))) | (~x15 & x18 & ~x19) | (x17 & (~x18 | (x15 & x18 & ~x19))))) : (~x13 & (x15 ? ((~x17 & (~x18 | (x18 & ~x19))) | (x17 & ((x05 & (x18 ^ x19)) | (~x18 & ~x19) | (~x05 & x18 & x19))) | (x05 & x18 & x19)) : ~x17)))) | (~x05 & (x12 ? (~x13 | (x13 & ~x16 & ((~x15 & (~x18 | (x17 & x18))) | (~x17 & (x18 | (x15 & ~x18)))))) : (x13 | (~x16 & ~x17 & ~x13 & ~x15)))) | (~x12 & ~x13 & (x15 ? ~x16 : x17)) | (x12 & x13 & x15 & ~x16 & x17))) | (~x05 & ~x12 & ~x13 & x15 & x16 & (x17 ? (x18 ^ x19) : (x18 & x19)))) : ~x05)))) | (~x14 & ((x02 & ~x03 & ~x04 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))) | (~x12 & x13 & ((x15 & ~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))))) | (x03 & ~x15 & x16 & x17 & x18 & x19 & (~x04 | (x04 & x05))))))))))))))));
  assign z28 = ~x08 & (x09 ? (~x10 | (x10 & x11)) : (x10 | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x10 & ~x11 & ~x14 & x15 & ~x16 & ~x17 & ~x36 & ~x37 & ~x38 & ~x39 & x40 & ((~x12 & x13 & x18) | (~x18 & ~x19 & x12 & ~x13)))));
  assign z29 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & (x10 | (~x10 & (x09 | (~x09 & ~x11 & (x36 | (~x36 & (x00 ? (~x01 & ~x02 & ~x14 & ((~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x12 & x13 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))))) : ((~x12 & x13 & ~x14 & ((x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))) | (x01 & (x15 ? (~x17 & ~x18 & ((x04 & ((((~x16 & x19) | (x05 & x16 & ~x19)) & (~x02 | (x02 & x03))) | (~x05 & x16 & (x03 ? ~x19 : ~x02)))) | (~x02 & ~x03 & ~x04) | ((~x16 ^ ~x19) & (x03 ? ~x04 : x02)))) : (x16 & x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))))) | (~x01 & ((~x14 & ((x02 & ~x03 & ~x04 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))) | (~x12 & x13 & ((x15 & ~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))))) | (x03 & ~x15 & x16 & x17 & x18 & x19 & (~x04 | (x04 & x05))))))) | (~x02 & ((~x03 & ~x04 & (x40 ? ((x14 & ((x16 & (x12 ? (x13 & ((x19 & (x05 ? (x17 ? x18 : ~x15) : (x18 & (~x15 | (x15 & x17))))) | (~x05 & ~x17 & (x15 | (~x15 & ~x18))) | (~x15 & x18 & ~x19) | (x17 & (~x18 | (x15 & x18 & ~x19))))) : (~x13 & (x15 ? ((~x17 & (~x18 | (x18 & ~x19))) | (x17 & ((x05 & (x18 ^ x19)) | (~x18 & ~x19) | (~x05 & x18 & x19))) | (x05 & x18 & x19)) : ~x17)))) | (~x05 & (x12 ? (~x13 | (x13 & ~x16 & ((~x15 & (~x18 | (x17 & x18))) | (~x17 & (x18 | (x15 & ~x18)))))) : (x13 | (~x16 & ~x17 & ~x13 & ~x15)))) | (~x12 & ~x13 & (x15 ? ~x16 : x17)) | (x12 & x13 & x15 & ~x16 & x17))) | (~x05 & ~x12 & ~x13 & x15 & x16 & (x17 ? (x18 ^ x19) : (x18 & x19)))) : ~x05)) | (~x14 & ((~x13 & ((~x03 & ~x04 & x40 & ((x16 & ((~x05 & ((~x15 & ((x12 & ~x19 & (x18 | (x17 & ~x18))) | (x17 & ~x18 & x19) | (~x17 & (~x18 | (x18 & x19))))) | (~x12 & (x17 ? (~x18 ^ x19) : (x18 ? ~x19 : x15))))) | (x12 & x15 & (~x17 | (x17 & (~x18 | (x18 & ~x19))))))) | (x17 & x18 & ((~x05 & ~x15 & (~x12 ^ x19)) | (x12 & x15 & x19))))) | (~x16 & ((~x03 & ~x04 & ~x05 & x40 & ((~x12 & ((x17 & (x15 ? x19 : ~x18)) | (~x15 & (x19 ? x18 : ~x17)))) | (~x17 & x19 & (x15 ^ ~x18)) | (x15 & ~x19 & (x18 | (x17 & ~x18))))) | (x12 & ((~x19 & ((~x15 & ((x17 & (x18 ? (x20 ? ((~x21 & (x03 ? (~x04 | (x04 & x27)) : x04)) | (~x03 & ~x04 & (x05 | (~x05 & x40)))) : (x21 & (x03 ? (x05 ? ((~x24 & (~x22 | (x22 & ~x23)) & (~x04 ^ x27)) | (~x04 & (x27 | (x22 & x23 & x24 & x25 & ~x27)))) : (~x04 | (x04 & x27 & (~x22 | (x22 & ~x24))))) : (x05 | (~x05 & (x04 | (~x04 & x40))))))) : (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05))))) | (~x03 & ~x04 & ~x05 & ~x18 & x40))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18 & x40 & (x38 | x39 | (~x38 & ~x39))))) | (~x03 & ((~x17 & x18 & x19 & x05 & x15) | (~x05 & ((~x17 & x18 & x40 & ~x04 & ~x15) | (x19 & ((~x17 & x18 & x04 & x15) | (~x04 & ~x18 & x40 & (x15 | (~x15 & x17 & x39))))))))))))))) | (~x03 & ~x04 & ~x05 & x12 & x13 & x40) | (~x12 & ((~x03 & ~x04 & ~x05 & x15 & ~x18 & x40 & ~x16 & ~x17) | (x13 & ((~x03 & ((~x15 & ((~x04 & ((x17 & ~x18 & ~x19 & x05 & x16) | (~x05 & ~x16 & x40))) | (x17 & x18 & x19 & x05 & x16))) | (~x04 & ~x05 & x16 & x40))) | (x18 & x19 & x16 & x17 & x04 & ~x05 & ~x15) | (x15 & ((~x17 & ~x18 & (x05 ? ~x03 : x04)) | (~x16 & ((x17 & (((~x19 | (~x18 & x19)) & (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05)))) | (~x05 & x40 & ~x03 & ~x04))) | (~x03 & ~x04 & ~x05 & ~x17 & x18 & x40 & (x38 | x39 | (~x38 & ~x39))))))))))))))))))))))))));
  assign z30 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & x19 & ~x36 & x40 & (~x17 | (x17 & (~x37 | x38 | ~x39 | (x37 & ~x38))));
  assign z33 = ~x08 & ~x09 & (x10 | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x10 & ~x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & x19 & ~x36 & x40 & (~x17 | (x17 & (~x37 | x38 | ~x39 | (x37 & ~x38))))));
  assign z34 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & ((x10 & (~x09 | (x09 & ~x11))) | (~x09 & ~x10 & ~x11 & (x36 | (~x36 & (x00 ? (~x01 & ~x02 & ~x14 & ((~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x12 & x13 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))))) : ((~x12 & x13 & ~x14 & ((x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))) | (x01 & (x15 ? (~x17 & ~x18 & ((x04 & ((((~x16 & x19) | (x05 & x16 & ~x19)) & (~x02 | (x02 & x03))) | (~x05 & x16 & (x03 ? ~x19 : ~x02)))) | (~x02 & ~x03 & ~x04) | ((~x16 ^ ~x19) & (x03 ? ~x04 : x02)))) : (x16 & x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))))) | (~x01 & ((~x14 & ((x02 & ~x03 & ~x04 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))) | (~x12 & x13 & ((x15 & ~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))))) | (x03 & ~x15 & x16 & x17 & x18 & x19 & (~x04 | (x04 & x05))))))) | (~x02 & ((~x03 & ~x04 & (x40 ? ((x14 & ((x16 & (x12 ? (x13 & ((x19 & (x05 ? (x17 ? x18 : ~x15) : (x18 & (~x15 | (x15 & x17))))) | (~x05 & ~x17 & (x15 | (~x15 & ~x18))) | (~x15 & x18 & ~x19) | (x17 & (~x18 | (x15 & x18 & ~x19))))) : (~x13 & (x15 ? ((~x17 & (~x18 | (x18 & ~x19))) | (x17 & ((x05 & (x18 ^ x19)) | (~x18 & ~x19) | (~x05 & x18 & x19))) | (x05 & x18 & x19)) : ~x17)))) | (~x05 & (x12 ? (~x13 | (x13 & ~x16 & ((~x15 & (~x18 | (x17 & x18))) | (~x17 & (x18 | (x15 & ~x18)))))) : (x13 | (~x16 & ~x17 & ~x13 & ~x15)))) | (~x12 & ~x13 & (x15 ? ~x16 : x17)) | (x12 & x13 & x15 & ~x16 & x17))) | (~x05 & ~x12 & ~x13 & x15 & x16 & (x17 ? (x18 ^ x19) : (x18 & x19)))) : ~x05)) | (~x14 & ((~x03 & ~x04 & ~x05 & x12 & x13 & x40) | (~x12 & ((~x03 & ~x04 & ~x05 & x15 & ~x18 & x40 & ~x16 & ~x17) | (x13 & ((~x03 & ((~x15 & ((~x04 & ((x17 & ~x18 & ~x19 & x05 & x16) | (~x05 & ~x16 & x40))) | (x17 & x18 & x19 & x05 & x16))) | (~x04 & ~x05 & x16 & x40))) | (x18 & x19 & x16 & x17 & x04 & ~x05 & ~x15) | (x15 & ((~x17 & ~x18 & (x05 ? ~x03 : x04)) | (~x16 & ((x17 & (((~x19 | (~x18 & x19)) & (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05)))) | (~x05 & x40 & ~x03 & ~x04))) | (~x03 & ~x04 & ~x05 & ~x17 & x18 & x40 & (x38 | x39 | (~x38 & ~x39))))))))))) | (~x13 & ((~x03 & ~x04 & x40 & ((x16 & ((~x05 & ((~x15 & ((x12 & ~x19 & (x18 | (x17 & ~x18))) | (x17 & ~x18 & x19) | (~x17 & (~x18 | (x18 & x19))))) | (~x12 & (x17 ? (~x18 ^ x19) : (x18 ? ~x19 : x15))))) | (x12 & x15 & (~x17 | (x17 & (~x18 | (x18 & ~x19))))))) | (x17 & x18 & ((~x05 & ~x15 & (~x12 ^ x19)) | (x12 & x15 & x19))))) | (~x16 & ((~x03 & ~x04 & ~x05 & x40 & ((~x12 & ((x17 & (x15 ? x19 : ~x18)) | (~x15 & (x19 ? x18 : ~x17)))) | (~x17 & x19 & (x15 ^ ~x18)) | (x15 & ~x19 & (x18 | (x17 & ~x18))))) | (x12 & ((~x03 & ((~x05 & ((x19 & ((~x04 & ~x18 & x40 & (x15 | (~x15 & x17))) | (~x17 & x18 & x04 & x15))) | (~x17 & x18 & x40 & ~x04 & ~x15))) | (~x17 & x18 & x19 & x05 & x15))) | (~x19 & ((~x15 & ((x17 & (x18 ? (x20 ? ((~x21 & (x03 ? (~x04 | (x04 & x27)) : x04)) | (~x03 & ~x04 & (x05 | (~x05 & x40)))) : (x21 & (x03 ? (x05 ? ((~x24 & (~x22 | (x22 & ~x23)) & (~x04 ^ x27)) | (~x04 & (x27 | (x22 & x23 & x24 & x25 & ~x27)))) : (~x04 | (x04 & x27 & (~x22 | (x22 & ~x24))))) : (x05 | (~x05 & (x04 | (~x04 & x40))))))) : (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05))))) | (~x03 & ~x04 & ~x05 & ~x18 & x40))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18 & x40 & (x38 | x39 | (~x38 & ~x39))))))))))))))))))))))));
  assign z35 = ~x08 & (x09 ? (~x10 | (x10 & x11)) : x10);
  assign z36 = ~x08 & (x09 ? (~x10 | (x10 & x11)) : (x10 | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x10 & ~x11 & x12 & ~x13 & ~x14 & ~x16 & ~x17 & ~x36 & x40 & ((~x15 & x18 & x19) | (x15 & ~x18 & ~x19 & ~x38 & ~x39)))));
  assign z37 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & ~x11 & (x09 ? x10 : (~x10 & (x36 | (~x36 & (x00 ? (~x01 & ~x02 & ~x14 & ((~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x12 & x13 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))))) : ((~x12 & x13 & ~x14 & ((x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))) | (x01 & (x15 ? (~x17 & ~x18 & ((x04 & ((((~x16 & x19) | (x05 & x16 & ~x19)) & (~x02 | (x02 & x03))) | (~x05 & x16 & (x03 ? ~x19 : ~x02)))) | (~x02 & ~x03 & ~x04) | ((~x16 ^ ~x19) & (x03 ? ~x04 : x02)))) : (x16 & x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))))) | (~x01 & ((~x14 & ((x02 & ~x03 & ~x04 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))) | (~x12 & x13 & ((x15 & ~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))))) | (x03 & ~x15 & x16 & x17 & x18 & x19 & (~x04 | (x04 & x05))))))) | (~x02 & ((~x03 & ~x04 & (x40 ? ((x14 & ((x16 & (x12 ? (x13 & ((x19 & (x05 ? (x17 ? x18 : ~x15) : (x18 & (~x15 | (x15 & x17))))) | (~x05 & ~x17 & (x15 | (~x15 & ~x18))) | (~x15 & x18 & ~x19) | (x17 & (~x18 | (x15 & x18 & ~x19))))) : (~x13 & (x15 ? ((~x17 & (~x18 | (x18 & ~x19))) | (x17 & ((x05 & (x18 ^ x19)) | (~x18 & ~x19) | (~x05 & x18 & x19))) | (x05 & x18 & x19)) : ~x17)))) | (~x05 & (x12 ? (~x13 | (x13 & ~x16 & ((~x15 & (~x18 | (x17 & x18))) | (~x17 & (x18 | (x15 & ~x18)))))) : (x13 | (~x16 & ~x17 & ~x13 & ~x15)))) | (~x12 & ~x13 & (x15 ? ~x16 : x17)) | (x12 & x13 & x15 & ~x16 & x17))) | (~x05 & ~x12 & ~x13 & x15 & x16 & (x17 ? (x18 ^ x19) : (x18 & x19)))) : ~x05)) | (~x14 & ((~x13 & ((~x03 & ~x04 & x40 & ((x16 & ((~x05 & ((~x15 & ((x12 & ~x19 & (x18 | (x17 & ~x18))) | (x17 & ~x18 & x19) | (~x17 & (~x18 | (x18 & x19))))) | (~x12 & (x17 ? (~x18 ^ x19) : (x18 ? ~x19 : x15))))) | (x12 & x15 & (~x17 | (x17 & (~x18 | (x18 & ~x19))))))) | (x17 & x18 & ((~x05 & ~x15 & (~x12 ^ x19)) | (x12 & x15 & x19))))) | (~x16 & ((~x03 & ~x04 & ~x05 & x40 & ((~x12 & ((x17 & (x15 ? x19 : ~x18)) | (~x15 & (x19 ? x18 : ~x17)))) | (~x17 & x19 & (x15 ^ ~x18)) | (x15 & ~x19 & (x18 | (x17 & ~x18))))) | (x12 & ((~x03 & ((~x05 & ((x19 & ((~x04 & ~x18 & x40 & (x15 | (~x15 & x17))) | (~x17 & x18 & x04 & x15))) | (~x17 & x18 & x40 & ~x04 & ~x15))) | (~x17 & x18 & x19 & x05 & x15))) | (~x19 & ((~x15 & ((x17 & (x18 ? (x20 ? ((~x21 & (x03 ? (~x04 | (x04 & x27)) : x04)) | (~x03 & ~x04 & (x05 | (~x05 & x40)))) : (x21 & (x03 ? (x05 ? ((~x24 & (~x22 | (x22 & ~x23)) & (~x04 ^ x27)) | (~x04 & (x27 | (x22 & x23 & x24 & x25 & ~x27)))) : (~x04 | (x04 & x27 & (~x22 | (x22 & ~x24))))) : (x05 | (~x05 & (x04 | (~x04 & x40))))))) : (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05))))) | (~x03 & ~x04 & ~x05 & ~x18 & x40))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18 & x40 & (x38 | x39 | (~x38 & ~x39))))))))))) | (~x03 & ~x04 & ~x05 & x12 & x13 & x40) | (~x12 & ((~x03 & ~x04 & ~x05 & x15 & ~x18 & x40 & ~x16 & ~x17) | (x13 & ((~x03 & ((~x15 & ((~x04 & ((x17 & ~x18 & ~x19 & x05 & x16) | (~x05 & ~x16 & x40))) | (x17 & x18 & x19 & x05 & x16))) | (~x04 & ~x05 & x16 & x40))) | (x18 & x19 & x16 & x17 & x04 & ~x05 & ~x15) | (x15 & ((~x17 & ~x18 & (x05 ? ~x03 : x04)) | (~x16 & ((x17 & (((~x19 | (~x18 & x19)) & (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05)))) | (~x05 & x40 & ~x03 & ~x04))) | (~x03 & ~x04 & ~x05 & ~x17 & x18 & x40 & (x38 | x39 | (~x37 & ~x38 & ~x39))))))))))))))))))))))));
  assign z38 = (~x02 & ~x03 & ~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x36) | (~x08 & ~x11 & (x09 ? x10 : (~x10 & (x36 | (~x36 & (x00 ? (~x01 & ~x02 & ~x14 & ((~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x12 & x13 & ((x16 & ((~x05 & ((x03 & ~x04 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x17 & ~x18 & ~x19 & ~x03 & x04 & x15))) | (~x03 & ((x18 & x19 & ~x15 & x17) | (~x17 & ~x18 & ~x19 & x05 & x15))))) | (~x03 & ~x04 & ~x05 & x15 & ~x17 & ~x18))))) : ((~x12 & x13 & ~x14 & ((x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))) | (x01 & (x15 ? (~x17 & ~x18 & ((x04 & ((((~x16 & x19) | (x05 & x16 & ~x19)) & (~x02 | (x02 & x03))) | (~x05 & x16 & (x03 ? ~x19 : ~x02)))) | (~x02 & ~x03 & ~x04) | ((~x16 ^ ~x19) & (x03 ? ~x04 : x02)))) : (x16 & x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))))) | (~x01 & ((~x14 & ((x02 & ~x03 & ~x04 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))) | (~x12 & x13 & ((x15 & ~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))))) | (x03 & ~x15 & x16 & x17 & x18 & x19 & (~x04 | (x04 & x05))))))) | (~x02 & ((~x03 & ~x04 & (x40 ? ((x14 & ((x16 & (x12 ? (x13 & ((x19 & (x05 ? (x17 ? x18 : ~x15) : (x18 & (~x15 | (x15 & x17))))) | (~x05 & ~x17 & (x15 | (~x15 & ~x18))) | (~x15 & x18 & ~x19) | (x17 & (~x18 | (x15 & x18 & ~x19))))) : (~x13 & (x15 ? ((~x17 & (~x18 | (x18 & ~x19))) | (x17 & ((x05 & (x18 ^ x19)) | (~x18 & ~x19) | (~x05 & x18 & x19))) | (x05 & x18 & x19)) : ~x17)))) | (~x05 & (x12 ? (~x13 | (x13 & ~x16 & ((~x15 & (~x18 | (x17 & x18))) | (~x17 & (x18 | (x15 & ~x18)))))) : (x13 | (~x16 & ~x17 & ~x13 & ~x15)))) | (~x12 & ~x13 & (x15 ? ~x16 : x17)) | (x12 & x13 & x15 & ~x16 & x17))) | (~x05 & ~x12 & ~x13 & x15 & x16 & (x17 ? (x18 ^ x19) : (x18 & x19)))) : ~x05)) | (~x14 & ((~x03 & ~x04 & ~x05 & x12 & x13 & x40) | (~x12 & ((~x03 & ~x04 & ~x05 & x15 & ~x18 & x40 & ~x16 & ~x17) | (x13 & ((~x03 & ((~x15 & ((~x04 & ((x17 & ~x18 & ~x19 & x05 & x16) | (~x05 & ~x16 & x40))) | (x17 & x18 & x19 & x05 & x16))) | (~x04 & ~x05 & x16 & x40))) | (x18 & x19 & x16 & x17 & x04 & ~x05 & ~x15) | (x15 & ((~x17 & ~x18 & (x05 ? ~x03 : x04)) | (~x16 & ((x17 & (((~x19 | (~x18 & x19)) & (x03 ? (~x04 & ~x05) : (x05 | (x04 & ~x05)))) | (~x05 & x40 & ~x03 & ~x04))) | (~x03 & ~x04 & ~x05 & ~x17 & x18 & x40 & (x38 | x39 | (~x37 & ~x38 & ~x39))))))))))) | (~x13 & ((~x03 & ~x04 & x40 & ((x16 & ((~x05 & ((~x15 & ((x12 & ~x19 & (x18 | (x17 & ~x18))) | (x17 & ~x18 & x19) | (~x17 & (~x18 | (x18 & x19))))) | (~x12 & (x17 ? (~x18 ^ x19) : (x18 ? ~x19 : x15))))) | (x12 & x15 & (~x17 | (x17 & (~x18 | (x18 & ~x19))))))) | (x17 & x18 & ((~x05 & ~x15 & (~x12 ^ x19)) | (x12 & x15 & x19))))) | (~x16 & ((~x03 & ~x04 & ~x05 & x40 & ((~x12 & ((x17 & (x15 ? x19 : ~x18)) | (~x15 & (x19 ? x18 : ~x17)))) | (~x17 & x19 & (x15 ^ ~x18)) | (x15 & ~x19 & (x18 | (x17 & ~x18))))) | (x12 & ((~x19 & ((~x04 & ((~x05 & ((~x15 & ((x17 & (x03 ? (~x18 | (x18 & ~x20 & x21)) : (x18 & x40 & (x20 | (~x20 & x21))))) | (~x03 & ~x18 & x40))) | (~x03 & x15 & ~x17 & ~x18 & x40 & (x38 | x39)))) | (~x15 & x17 & x18 & ((x20 & (x03 ? ~x21 : x05)) | (x03 & x05 & ~x20 & x21 & (x27 | (~x27 & (x22 ? (x23 ? (x24 & x25) : ~x24) : ~x24)))))))) | (~x15 & x17 & (x03 ? (x04 & x18 & x27 & (x20 ? ~x21 : (x21 & ((~x05 & ~x22) | (~x24 & (x05 ? (~x22 | (x22 & ~x23)) : x22)))))) : (((x05 | (x04 & ~x05)) & (~x18 | (x18 & ~x20 & x21))) | (x20 & ~x21 & x04 & x18)))))) | (~x03 & x19 & ((~x05 & ((~x04 & ~x18 & x40 & (x15 | (~x15 & x17))) | (~x17 & x18 & x04 & x15))) | (~x17 & x18 & x05 & x15))))))))))))))))))))));
  assign z40 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x13 & ~x14 & ~x16 & ~x17 & ~x36 & x40 & ((x15 & ~x18 & ~x19 & ~x38 & ~x39) | (~x15 & x18));
  assign z41 = ~x01 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x14 & ((~x04 & ((~x02 & ((~x05 & ((x13 & ((~x12 & ((x16 & (x00 ? (x03 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) : (~x03 & ~x15 & x40 & (x19 ? ~x18 : ~x17)))) | (~x00 & x15 & ~x16 & x17 & ((x03 & ~x19) | (x19 & x40 & ~x03 & x18))))) | (~x00 & ~x03 & x12 & x28 & x40 & (x15 | (~x15 & x24 & x25 & x26))))) | (~x00 & x12 & ~x13 & x17 & ((~x03 & x40 & (x18 ^ x19) & (x15 ^ x16)) | (x03 & ~x15 & ~x16 & x18 & ~x19 & ~x20 & x21 & x22 & ~x23 & x24 & ~x27))))) | (~x00 & x03 & x05 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & (x20 ? (~x21 & ~x27) : (x21 & (x22 ? ((~x23 & (x24 ^ ~x27)) | (x23 & x24 & ~x26 & x27)) : (~x24 & ~x27))))))) | (~x00 & x02 & ~x03 & x12 & ~x13 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x05 ? (x20 & ~x21) : (~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))))) | (~x00 & ~x02 & x04 & x05 & x12 & ~x13 & ~x16 & x18 & ((~x17 & x19 & ~x03 & x15) | (x21 & x22 & ~x23 & ~x24 & x27 & x03 & ~x15 & x17 & ~x19 & ~x20))))) | (~x04 & ~x05 & x12 & ~x00 & ~x02 & ~x03 & x13 & x14 & x15 & x16 & ~x17 & x40));
  assign z42 = ~x00 & ~x01 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x04 & ((x12 & ((~x13 & ((~x14 & ((~x16 & ((x17 & ((~x15 & x18 & ~x19 & ((~x20 & x21 & ((~x24 & ((x02 & ~x03 & ~x05 & x27 & (~x22 | (x22 & ~x23))) | (~x02 & x03 & x05 & x22 & ~x23 & ~x27))) | (~x02 & x03 & x05 & x22 & ~x23 & x24 & x27))) | (x20 & ~x21 & x27 & x02 & ~x03 & x05))) | (~x02 & ~x03 & ~x05 & x19 & x40 & x15 & ~x18))) | (~x02 & ~x03 & ~x05 & ~x19 & x40 & x15 & x18))) | (~x02 & ~x03 & ~x05 & ~x15 & ~x18 & x19 & x40 & x16 & x17))) | (~x02 & ~x03 & ~x05 & x14 & x15 & x40))) | (~x02 & ~x03 & ~x05 & x13 & ~x14 & x30 & x32 & x33 & x34 & x40))) | (~x02 & ~x03 & ~x05 & ~x12 & x13 & x14 & x15 & x40))) | (x17 & x18 & ~x19 & ~x20 & x21 & x22 & ~x23 & ~x24 & x27 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x04 & x05 & ~x02 & x03));
  assign z43 = ~x01 & ~x02 & ~x04 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x00 & ((x12 & ((x17 & (x05 ? ((~x03 & x40 & ((x13 & x14 & (x16 ? ~x18 : x15)) | (x15 & x16 & ~x18 & ~x13 & ~x14))) | (x18 & ((~x03 & x13 & x14 & x16 & x40 & (x19 | (x15 & ~x19))) | (~x13 & ~x14 & ((x19 & x40 & ~x03 & x15) | (~x19 & ((x16 & x40 & ~x03 & x15) | (x03 & ~x15 & ~x16 & ~x20 & x21 & x22 & x23 & x24 & (x27 ? x26 : x25))))))))) : (~x15 & ((~x03 & x40 & (x13 ? (x14 & ~x16 & (x18 ^ x19)) : (~x14 & x16 & ~x18 & ~x19 & (~x38 | ~x39)))) | (~x16 & ~x18 & ~x19 & x03 & ~x13 & ~x14))))) | (~x03 & x40 & (x13 ? (~x15 & ((x05 & x14 & x16 & (x19 ? ~x17 : x18)) | (~x05 & ~x14 & x20 & x21 & x22 & x23 & x29))) : ((~x14 & ~x17 & (x05 ? (x15 & x16) : ((~x15 & x16 & x18) | (~x18 & x19 & x15 & ~x16)))) | (~x05 & x14 & ~x15)))))) | (~x03 & ~x12 & x40 & ((~x15 & ((x14 & (x05 ? (~x13 & x17) : (x13 | (~x13 & ~x16 & ~x17 & x18 & x19)))) | (~x05 & x13 & ~x14 & (~x16 | (x18 & x19 & x16 & ~x17))))) | (x05 & ~x13 & x14 & ((x16 & ~x17) | (x15 & (~x16 | (x16 & x17))))))))) | (x17 & ~x18 & ~x19 & ~x14 & ~x15 & ~x16 & ~x05 & x12 & ~x13 & x00 & ~x03));
  assign z44 = ~x00 & ~x01 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & ~x36 & (x02 ? (~x03 & ~x04 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))) : (x04 ? (x27 & ((~x03 & x20 & ~x21) | (~x20 & x21 & ((~x24 & (((~x22 | (x22 & ~x23)) & (~x03 | (x03 & x05))) | (x03 & ~x05 & x22 & x23))) | (x03 & ~x05 & ~x22 & x24))))) : ((x05 & (x20 ? (~x21 & (~x03 | (x03 & ~x27))) : (x21 & (((~x22 | (x22 & ~x23)) & (x27 ? (~x03 | (x03 & x24)) : ~x24)) | (x22 & x23 & (x24 ? ((~x26 & x27) | (x03 & x25 & ~x27)) : x27)))))) | (~x05 & ((~x20 & x21 & (x03 ? (~x27 & (x24 | (x22 & x23 & ~x24))) : x40)) | (~x03 & x20 & x40))) | (x21 & x22 & x03 & ~x20 & x23 & x24 & x26 & x27))));
  assign z45 = ~x01 & ~x02 & ~x04 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((x17 & ~x18 & ~x19 & ~x14 & ~x15 & ~x16 & ~x05 & x12 & ~x13 & x00 & ~x03) | (~x00 & ((~x03 & ((x12 & ((~x13 & ((~x14 & ((x17 & ((~x19 & (x05 ? (~x15 & ~x16 & x18 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : (x40 & ((x15 & (~x16 | (x16 & ~x18))) | (x18 & (x16 | (~x15 & ~x16 & (x20 | (~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))))))))) | (~x05 & x19 & x40 & (x18 | (x16 & ~x18))))) | (~x05 & x40 & ((~x18 & (x15 ? (x16 ? ~x17 : x19) : (~x16 & ~x19))) | (x16 & ~x17 & x18 & (x19 | (x15 & ~x19))))))) | (~x05 & x14 & x40))) | (~x05 & x13 & x14 & x40 & ((x17 & ((x15 & (x16 ? (x18 & ~x19) : ~x18)) | (~x16 & x18) | (x16 & (~x18 | (x18 & x19))))) | (x15 & ~x17) | (~x15 & ((x16 & (x19 ? ~x17 : x18)) | (~x18 & (x19 ? ~x16 : ~x17)))))))) | (~x05 & ~x12 & ~x13 & x14 & x40 & ((~x16 & (x15 | (~x15 & x18 & x19))) | (x16 & ~x17) | (x17 & (((~x18 | (x18 & ~x19)) & (~x15 | (x15 & x16))) | (x16 & x18 & x19))))))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & x03 & ~x05 & x12 & ~x13 & ~x14))));
  assign z46 = ~x00 & ~x01 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x04 & ((x12 & ((x17 & (x02 ? (~x03 & ~x13 & ~x14 & ~x15 & ~x16 & x18 & ~x19 & x27 & ((x20 & ~x21) | (~x05 & ~x20 & x21 & ~x24 & (~x22 | (x22 & ~x23))))) : ((x18 & ((~x05 & ((~x13 & ~x14 & ((x19 & x40 & ~x03 & x15) | (~x19 & ((x16 & x40 & ~x03 & x15) | (~x15 & ~x16 & x21 & (x03 ? (~x20 & ~x27 & (x24 | (x22 & x23 & ~x24))) : (x20 & x40))))))) | (~x03 & x13 & x14 & x40 & (~x16 | (x16 & (x19 | (x15 & ~x19))))))) | (x03 & ~x13 & ~x14 & ~x15 & ~x16 & ~x19 & ((x05 & (x20 ? (~x21 & ~x27) : (x21 & (((~x22 | (x22 & ~x23)) & (x24 ^ ~x27)) | (x22 & x23 & (x24 ? (x27 ? ~x26 : x25) : x27)))))) | (~x20 & x21 & x22 & x23 & x24 & x26 & x27))))) | (~x03 & ~x05 & ~x18 & x40 & ((x13 & x14 & (x16 | (x15 & ~x16))) | (x15 & x16 & ~x13 & ~x14)))))) | (~x02 & ~x03 & ~x05 & x40 & ((x13 & x14 & ~x15 & ((x16 & (x19 ? ~x17 : x18)) | (~x18 & (x19 ? ~x16 : ~x17)))) | (~x13 & ~x14 & x15 & x16 & ~x17))))) | (~x02 & ~x03 & ~x05 & ~x12 & ~x13 & x14 & x40 & ((~x16 & (x15 | (~x15 & x18 & x19))) | (x16 & ~x17) | (x17 & (((~x18 | (x18 & ~x19)) & (~x15 | (x15 & x16))) | (x16 & x18 & x19))))))) | (~x02 & x03 & x04 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & ~x20 & x21 & x27 & ((~x24 & (x05 ? (~x22 | (x22 & ~x23)) : (x22 & x23))) | (~x05 & ~x22 & x24))));
  assign z47 = ~x08 & ((~x10 & (x09 | (~x00 & ~x01 & ~x09 & ~x11 & ~x36 & ((~x03 & ((~x04 & ((~x13 & ((x17 & ((x12 & ~x14 & ((~x19 & ((~x15 & ((~x02 & ~x05 & x16 & ~x18 & x40 & (~x38 | ~x39)) | (~x16 & x18 & ((x27 & (x02 ? ((x05 & x20 & ~x21) | (~x05 & ~x20 & x21 & ~x22 & ~x24)) : (~x05 & x40 & (x20 ? ~x21 : (x21 & (~x22 | (x22 & (~x23 | (x23 & (~x24 | (x24 & ~x26))))))))))) | (~x02 & ~x05 & x20 & x21 & x40))))) | (~x02 & ~x05 & x15 & x16 & x18 & x40))) | (~x02 & ~x05 & x15 & x40 & (x18 ? x19 : x16)))) | (~x02 & ~x05 & ~x12 & x14 & x40 & (((~x18 | (x18 & ~x19)) & (~x15 | (x15 & x16))) | (x16 & x18 & x19))))) | (~x02 & ~x05 & x40 & ((x15 & (x12 ? (~x14 & ~x17 & (x16 | (~x37 & ~x38 & ~x39 & ~x16 & ~x18 & ~x19))) : (x14 & ~x16))) | (~x12 & x14 & ((x16 & ~x17) | (x18 & x19 & ~x15 & ~x16))))))) | (~x02 & ~x05 & x13 & x40 & ((x12 & x14 & ((x15 & ~x16 & x17) | (x16 & ((~x15 & (x19 ? ~x17 : x18)) | (x17 & (~x18 | (x18 & x19))) | (x15 & (~x17 | (x17 & x18 & ~x19))))))) | (x15 & ~x16 & ~x12 & ~x14 & ~x37 & ~x38 & ~x39 & ~x17 & x18))))) | (~x02 & x04 & ~x05 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))))) | (~x02 & x03 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & ~x20 & x21 & ((x27 & ((x04 & ~x05 & (x22 ? (x23 & ~x24) : x24)) | (~x04 & x05 & x22 & x23 & x24 & x26))) | (~x04 & x05 & x22 & x25 & ~x27 & x23 & x24))))))) | (x09 & x10 & x11));
  assign z48 = ~x01 & ~x02 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x00 & ((~x03 & x40 & ((~x13 & (((~x18 | (x18 & ~x19)) & ((~x12 & x14 & x17 & (~x15 | (x15 & x16))) | (x15 & x16 & ~x17 & x12 & ~x14))) | (x16 & (x12 ? (~x14 & (x17 ? (x18 ? ~x19 : (x19 | (~x19 & (x15 | (~x15 & (~x38 | ~x39)))))) : (x18 & x19))) : (x14 & (~x17 | (x17 & x18 & x19))))) | (~x16 & (x12 ? (~x14 & (x15 ? (x19 ? ~x18 : x17) : (~x18 & ~x19))) : (x14 & (x15 | (~x15 & x18 & x19))))) | (x12 & (x14 | (x18 & x19 & ~x14 & x17))))) | (x12 & x13 & x14 & ((x17 & ((x15 & (~x16 | (x16 & x18 & ~x19))) | (x16 & (~x18 | (x18 & x19))) | (~x15 & x18 & ~x19))) | (x15 & ~x17) | (~x15 & ((~x16 & ~x18 & x19) | (~x17 & (x16 ? (x19 | (x18 & ~x19)) : (~x18 & ~x19))))))))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & ~x13 & ~x14 & x03 & x12))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & x00 & ~x03 & x12 & ~x13 & ~x14));
  assign z49 = ~x08 & ~x09 & ~x10 & ~x11 & ~x12 & x13 & ~x14 & ~x36 & (x00 ? (~x01 & ~x02 & ~x03 & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18 & ((x16 & ~x19) | (~x16 & x19 & ~x04 & ~x05))))) : ((x02 & ~x15 & x16 & x17 & x18 & x19 & (~x03 | (x03 & x04 & ~x05))) | (x01 & (x15 ? (~x17 & ~x18 & ((x04 & ((((~x16 & x19) | (x05 & x16 & ~x19)) & (~x02 | (x02 & x03))) | (~x05 & x16 & (x03 ? ~x19 : ~x02)))) | (~x02 & ~x03 & ~x04) | ((~x16 ^ ~x19) & (x03 ? ~x04 : x02)))) : (x16 & x17 & x18 & x19 & (~x02 | (x02 & x03 & (~x04 | (x04 & x05))))))) | (~x01 & (x15 ? (~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05))) | (~x02 & ((x04 & ~x05) | (~x03 & (x05 | (~x04 & ~x05 & x40))))))) : (x16 & x17 & x18 & x19 & ((x03 & (~x04 | (x04 & x05))) | (~x02 & ((x04 & ~x05) | (~x03 & (x05 | (~x04 & ~x05 & x40)))))))))));
  assign z50 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & (x00 ? (~x01 & ~x02 & ~x03 & ~x14 & ((~x12 & x13 & ((x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17)) & (~x04 | (x04 & ~x05))) | (~x18 & x19 & ~x16 & ~x17 & ~x04 & ~x05 & x15))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & ~x04 & ~x05 & x12 & ~x13))) : ((x13 & ((~x01 & ((~x02 & ((~x03 & ~x04 & ~x05 & x40 & ((x12 & (~x14 | (x14 & ((x15 & ~x17) | (~x15 & ~x16 & x17 & ~x18 & x19))))) | (~x12 & ~x14 & ~x15 & ~x18 & x19 & x16 & ~x17))) | (x04 & ~x12 & ~x14 & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18 & (~x16 ^ ~x19)))))) | (x03 & ~x04 & ~x12 & ~x14 & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18 & (~x16 ^ ~x19)))))) | (~x12 & ~x14 & ((x17 & x18 & x19 & ~x15 & x16) | (x15 & ~x17 & ~x18 & (~x16 ^ ~x19))) & ((x02 & (~x03 | (x03 & x04))) | (x01 & (~x02 | (x02 & x03 & ~x04))))))) | (~x01 & ~x02 & ~x04 & x12 & ~x13 & ((~x16 & x17 & ~x18 & ~x19 & ~x14 & ~x15 & x03 & ~x05) | (~x03 & ((x05 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ~x19) | (~x05 & x40 & (x14 | (~x14 & ((~x15 & x17 & ((x18 & x19) | (x16 & (x18 ^ x19)))) | (~x16 & ((~x18 & ~x19 & ~x15 & x17) | (x15 & ((~x18 & x19) | (x17 & x18 & ~x19)))))))))))))));
  assign z51 = ~x02 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x03 & (x00 ? (~x01 & ~x14 & ((~x15 & ~x16 & x17 & ~x18 & ~x19 & ~x04 & ~x05 & x12 & ~x13) | (x04 & ~x12 & x13 & x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))))) : ((~x14 & ((x13 & ((~x12 & ((~x17 & ~x18 & ((x15 & (x01 ? ((x04 & ~x05 & x16 & x19) | (~x16 & ~x19 & ~x04 & x05)) : (~x04 & ((x05 & (~x16 ^ ~x19)) | (x19 & x40 & ~x05 & ~x16))))) | (~x01 & ~x04 & ~x05 & x16 & x40 & (~x19 | (~x15 & x19))))) | (~x01 & ~x04 & x17 & x18 & x19 & (x05 ? (~x15 & x16) : (x40 & (x15 ^ x16)))))) | (~x01 & ~x04 & ~x05 & x12 & x40 & (x15 | (~x17 & ~x18 & ~x19 & ~x15 & x16))))) | (~x01 & ~x04 & x12 & ~x13 & ((~x05 & x40 & ((~x16 & (x15 ? (x19 ? ~x18 : x17) : (~x18 & ~x19))) | (~x15 & x17 & ((x18 & x19) | (x16 & (x18 ^ x19)))))) | (x17 & ~x18 & ~x19 & x05 & ~x15 & ~x16))))) | (~x01 & ~x04 & ~x05 & x12 & x14 & x40 & (~x13 | (x13 & (x15 ? ~x17 : ((~x17 & ~x18 & ~x19) | (~x16 & x17 & x19))))))))) | (~x01 & x03 & ~x04 & ~x05 & ~x14 & ((x00 & ~x12 & x13 & x16 & ((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17))) | (~x16 & x17 & ~x18 & ~x19 & ~x13 & ~x15 & ~x00 & x12))));
  assign z52 = ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x14 & ((~x01 & ((~x12 & x13 & ((~x02 & ((~x04 & ((x16 & ((((x18 & x19 & ~x15 & x17) | (~x18 & ~x19 & x15 & ~x17)) & ((~x03 & x05) | (x00 & x03 & ~x05))) | (~x05 & ~x15 & ~x00 & ~x03 & ~x19 & x40 & ~x17 & ~x18))) | (~x00 & ~x03 & x15 & ~x16 & x19 & ((x05 & ~x17 & ~x18) | (x18 & x40 & ~x05 & x17))))) | (~x00 & x15 & ~x17 & ~x18 & (x05 ? ~x03 : x04) & (~x16 ^ x19)))) | (~x00 & x15 & ~x17 & ~x18 & ((x02 & (~x03 | (x03 & x04 & ~x05))) | (x03 & (~x04 | (x04 & x05)))) & (~x16 ^ x19)))) | (~x00 & ~x02 & ~x03 & ~x04 & ~x05 & x12 & ~x13 & ~x16 & ~x18 & ~x19 & x40 & (~x15 ^ x17)))) | (~x00 & x01 & ~x02 & ~x03 & ~x04 & ~x12 & x13 & x15 & ~x17 & ~x18 & ((x16 & x19) | (~x05 & ~x16 & ~x19))))) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x12 & ~x19 & x40 & ~x17 & ~x18 & ~x15 & ~x16 & x13 & x14));
  assign z53 = ~x02 & ~x03 & ~x04 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x00 & ((~x01 & ((~x14 & ((~x18 & ((~x19 & (x05 ? ((x12 & ~x13 & ~x15 & ~x16 & x17) | (~x12 & x13 & x15 & x16 & ~x17)) : (x15 & x40 & ((~x16 & x17 & x12 & ~x13) | (~x12 & x13 & x16 & ~x17))))) | (~x05 & ~x12 & x13 & ~x17 & x19 & x40 & (x15 | (~x15 & x16))))) | (~x05 & x13 & x40 & (x12 ? x15 : (x17 & x18 & x19 & (x15 ^ x16)))))) | (~x05 & x12 & x13 & x14 & x40 & (x15 ? (x16 & ~x17) : ((x18 & x19 & ~x16 & x17) | (~x18 & ~x19 & x16 & ~x17)))))) | (x01 & x05 & ~x12 & x13 & ~x14 & x15 & x16 & ~x17 & ~x18 & x19))) | (x00 & ~x01 & x05 & ~x12 & x13 & x17 & x18 & x19 & ~x14 & ~x15 & x16));
  assign z54 = ~x00 & ~x01 & ~x02 & ~x03 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x05 & ((~x14 & ((x13 & ((~x12 & ((x19 & ((x04 & ((~x15 & x16 & x17 & x18) | (x15 & ~x16 & ~x17 & ~x18))) | (~x04 & x15 & ~x16 & x17 & x18 & x40))) | (~x17 & ~x18 & x40 & ~x04 & ~x15 & x16))) | (~x04 & x12 & x40 & (x15 | (~x15 & ((x17 & x18) | (~x18 & x19 & x16 & ~x17))))))) | (~x04 & x12 & ~x13 & ~x16 & ~x18 & ~x19 & x40 & (~x15 ^ x17)))) | (~x04 & x12 & x13 & x14 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & x40))) | (~x04 & x05 & ~x12 & x13 & ~x14 & ~x17 & ~x18 & ~x19 & x15 & x16));
  assign z55 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & x13 & x15 & ~x36 & x40 & (~x14 | (x14 & x16 & ~x17 & (x18 ^ x19)));
  assign z56 = ~x00 & ~x01 & ~x02 & ~x03 & ~x08 & ~x09 & ~x10 & ~x11 & x13 & ~x14 & ~x36 & ((~x05 & (x04 ? (~x12 & x19 & ((~x15 & x16 & x17 & x18) | (x15 & ~x16 & ~x17 & ~x18))) : (x12 & x40 & (x15 | (~x15 & x16 & x17 & x18))))) | (~x18 & ~x19 & x16 & ~x17 & ~x04 & x05 & ~x12 & x15));
  assign z57 = ~x00 & ~x01 & ~x02 & ~x03 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((x13 & ((~x05 & ((~x14 & ((~x12 & ((x19 & ((x04 & ((~x15 & x16 & x17 & x18) | (x15 & ~x16 & ~x17 & ~x18))) | (~x17 & ~x18 & x40 & ~x04 & x16))) | (~x19 & x40 & ~x17 & ~x18 & ~x04 & x15 & ~x16))) | (~x04 & x12 & x40 & (x15 | (~x15 & x16 & ~x17 & ~x18 & x19))))) | (~x04 & x12 & x14 & ~x17 & x40 & x15 & x16))) | (~x17 & ~x18 & ~x19 & x15 & x16 & ~x04 & x05 & ~x12 & ~x14))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & ~x04 & x05 & x12 & ~x13 & ~x14));
  assign z58 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x08 & ~x09 & ~x10 & ~x11 & ~x14 & ~x18 & ~x36 & ((~x05 & ~x12 & x13 & x15 & ~x17 & x40 & (~x16 ^ x19)) | (x05 & x12 & ~x13 & x17 & ~x19 & ~x15 & ~x16));
  assign z59 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & x13 & x15 & ~x36 & x40 & (~x14 | (x14 & x16 & ~x17));
  assign z60 = ~x36 & ~x19 & ~x18 & x17 & x16 & ~x15 & ~x14 & x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z61 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x14 & x15 & ~x16 & ~x17 & ~x36 & ~x37 & ~x38 & ~x39 & x40 & ((~x12 & x13 & x18) | (~x18 & ~x19 & x12 & ~x13));
  assign z62 = ~x00 & ~x01 & ~x02 & ~x04 & ~x09 & ~x36 & ((~x03 & (x08 ? ~x05 : (~x10 & ~x11 & x40 & ((x16 & (x05 ? ((x14 & (x12 ? (x13 & ((~x15 & (x19 ? ~x17 : x18)) | (x17 & (~x18 | (x18 & (x19 | (x15 & ~x19))))))) : (~x13 & (~x17 | (x15 & x17))))) | (x12 & ~x13 & ~x14 & x15 & (~x17 | (x17 & (~x18 | (x18 & ~x19)))))) : (~x12 & ~x14 & ((x15 & (x18 ? ((x17 & x19) | (x13 & (~x17 | (x17 & ~x19)))) : x17)) | (~x13 & (~x17 | (x17 & x18 & ~x19))))))) | (~x16 & ((x14 & ((x05 & x15 & (x12 ? (x13 & x17) : ~x13)) | (~x18 & ~x19 & ~x15 & x17 & ~x05 & x12 & x13))) | (~x05 & ~x13 & ((~x12 & (x15 ? ~x14 : ((~x17 & ~x18 & ~x19) | (~x14 & (x19 ? ~x17 : x18))))) | (~x15 & x17 & x12 & ~x14 & ~x18 & x19 & x37 & ~x38))))) | (~x13 & x17 & (x05 ? ((~x12 & x14 & ~x15) | (x12 & ~x14 & x15 & x18 & x19)) : (~x12 & ~x14 & ~x15 & (~x18 | (x18 & x19))))))))) | (x03 & ~x05 & ~x08 & ~x10 & ~x11 & ~x12 & ~x16 & x17 & ~x18 & x13 & ~x14 & x15));
  assign z63 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x09 & ~x36 & (x08 | (~x08 & ~x10 & ~x11 & ~x14 & ~x16 & x37 & ~x38 & x40 & ((x12 & ~x13 & ~x18 & ((~x15 & x17 & x19) | (x15 & ~x17 & ~x19 & ~x39))) | (~x12 & x13 & x15 & ~x17 & x18 & ~x39))));
  assign z64 = x40 & ~x39 & ~x38 & ~x37 & ~x36 & x19 & x18 & ~x17 & ~x16 & x15 & ~x14 & x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x05 & ~x04 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z65 = ~x01 & ~x02 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x15 & ~x16 & x17 & ~x18 & ~x19 & x00 & ~x03 & x12 & ~x13 & ~x14) | (~x00 & ((~x15 & ~x16 & x17 & ~x18 & ~x19 & ~x13 & ~x14 & x03 & x12) | (~x03 & x40 & ((x12 & (x13 ? ((x14 & ~x16 & ((x15 & ~x17) | (~x18 & x19 & ~x15 & x17))) | (~x17 & ~x18 & ~x19 & ~x14 & ~x15 & x16)) : (x14 | (~x14 & ((~x15 & x17 & ((x18 & x19) | (x16 & (x18 ^ x19)))) | (~x16 & ((~x18 & ~x19 & ~x15 & x17) | (x15 & ((~x18 & x19) | (x17 & x18 & ~x19)))))))))) | (~x12 & x13 & ~x14 & x15 & ~x16 & x17 & ~x18 & x19))))));
  assign z66 = ~x00 & ~x01 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x13 & ~x14 & ~x15 & x17 & ~x36 & ((~x02 & ((~x03 & (x04 ? (~x16 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : (x05 ? (~x16 & x18 & ~x19 & (x20 ? ~x21 : (x21 & (((x27 | (~x24 & ~x27)) & (~x22 | (x22 & ~x23))) | (x22 & x23 & x27 & (~x24 | (x24 & ~x26))))))) : (x40 & ((x19 & (x16 ^ x18)) | (~x16 & x18 & ~x19 & (x20 | (~x20 & x21)))))))) | (x03 & ~x04 & x05 & ~x16 & x18 & ~x19 & x20 & ~x21 & ~x27))) | (x18 & ~x19 & x20 & ~x21 & x27 & x02 & ~x03 & ~x04 & ~x16));
  assign z67 = ~x00 & ~x01 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x19 & ~x36 & ((x18 & ~x20 & x21 & (((~x22 | (x22 & ~x23)) & ((~x02 & x03 & x05 & (x04 ? (~x24 & x27) : (x24 ^ ~x27))) | (x02 & ~x03 & ~x04 & ~x05 & ~x24 & x27))) | (~x02 & x03 & ((x27 & (x04 ? (~x05 & (x22 ? (x23 & ~x24) : x24)) : (x22 & x23 & ((x24 & x26) | (x05 & (~x24 | (x24 & ~x26))))))) | (~x04 & ~x27 & ((~x05 & (x24 | (x22 & x23 & ~x24))) | (x23 & x24 & x25 & x05 & x22))))))) | (~x02 & ~x03 & ~x04 & ~x05 & ~x18 & x40));
  assign z68 = ~x01 & ~x02 & ~x03 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x36 & ((~x00 & (x04 ? (~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & x27 & (x20 ? ~x21 : (x21 & ~x24 & (~x22 | (x22 & ~x23))))) : (x05 ? (~x13 & ~x14 & ~x15 & ~x16 & x17 & x18 & ~x19 & (x20 ? ~x21 : (x21 & (((x27 | (~x24 & ~x27)) & (~x22 | (x22 & ~x23))) | (x22 & x23 & x27 & (~x24 | (x24 & ~x26))))))) : (x40 & ((x15 & ((x14 & (~x13 | (~x17 & x18 & x13 & ~x16))) | (~x13 & ~x14 & ~x16 & x17 & (x18 ^ x19)))) | (~x13 & ~x14 & ~x15 & x17 & (x16 ? (x18 ^ x19) : (x18 & ~x19 & (x20 | (~x20 & x21)))))))))) | (~x15 & ~x16 & x17 & ~x18 & ~x19 & x00 & ~x04 & ~x05 & ~x13 & ~x14));
  assign z69 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & x13 & x15 & ~x36 & x40 & ((~x14 & ~x16) | (~x17 & ~x19 & x14 & x16));
  assign z70 = ~x00 & ~x01 & ~x02 & ~x04 & ~x08 & ~x09 & ~x10 & ~x11 & ~x36 & ((~x03 & x40 & ((~x16 & ((x14 & ((x05 & x15 & (x12 ? (x13 & x17) : ~x13)) | (~x18 & ~x19 & ~x15 & x17 & ~x05 & x12 & x13))) | (~x05 & ~x13 & ((~x12 & (x15 ? ~x14 : ((~x17 & ~x18 & ~x19) | (~x14 & (x19 ? ~x17 : x18))))) | (~x15 & x17 & x12 & ~x14 & ~x18 & x19 & x37 & ~x38))))) | (~x13 & x17 & (x05 ? ((~x12 & x14 & ~x15) | (x12 & ~x14 & x15 & x18 & x19)) : (~x12 & ~x14 & ~x15 & (~x18 | (x18 & x19))))) | (x16 & (x05 ? ((x14 & (x12 ? (x13 & ((~x15 & (x19 ? ~x17 : x18)) | (x17 & (~x18 | (x18 & (x19 | (x15 & ~x19))))))) : (~x13 & (~x17 | (x15 & x17))))) | (x12 & ~x13 & ~x14 & x15 & (~x17 | (x17 & (~x18 | (x18 & ~x19)))))) : ((x15 & ((x13 & (x12 ? (~x14 | (x14 & ~x17 & x19)) : (~x14 & x18 & (~x17 | (x17 & ~x19))))) | (~x12 & ~x14 & x17 & (~x18 | (x18 & x19))))) | (~x12 & ~x13 & ~x14 & (~x17 | (x17 & x18 & ~x19)))))))) | (x03 & ~x05 & ~x12 & x13 & ~x16 & x17 & ~x18 & ~x14 & x15));
  assign z71 = ~x10 & ~x08 & x09;
  assign z72 = ~x08 & ~x11 & (x09 ? x10 : (~x10 & (x36 | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x36 & (~x40 | (~x14 & x40 & (((x38 | x39) & ((x12 & ~x13 & ~x18 & ~x19 & (x15 ? (~x16 & ~x17) : (x16 & x17))) | (~x16 & ~x17 & x18 & ~x12 & x13 & x15))) | (x12 & ~x13 & ~x15 & ~x16 & x17 & ~x18 & x19 & x39))))))));
  assign z01 = 1'b0;
  assign z31 = 1'b0;
  assign z32 = 1'b0;
  assign z39 = 1'b0;
endmodule