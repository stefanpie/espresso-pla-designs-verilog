module pla__test2 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34;
  assign z00 = (~x09 & ((x03 & ((~x10 & (x04 ? ((x08 & ((((x01 & x02 & x05 & x07) | (~x01 & ~x02 & ~x05 & ~x07)) & (x00 ^ x06)) | (~x00 & ~x05 & ~x06 & (x01 ? (~x02 & x07) : (x02 & ~x07))))) | (~x05 & x06 & x07 & ~x08 & (x00 ? (x01 & ~x02) : (~x01 & x02)))) : ((x05 & ((x06 & ((~x07 & (x00 ? (x01 ? (~x02 & ~x08) : x08) : (~x02 & ~x08))) | (~x00 & x02 & x07 & (x01 ^ x08)))) | (~x00 & x01 & ~x02 & ~x06 & x07 & x08))) | (x00 & ~x01 & ~x02 & ~x05 & ~x06 & ~x07 & ~x08)))) | (x10 & ((x06 & (x01 ? (~x04 & ((x00 & ((x02 & x08 & (~x07 | (x05 & x07))) | (~x02 & ~x05 & x07 & ~x08))) | (~x00 & ~x02 & ~x05 & x08))) : (x04 & ((~x08 & ((~x00 & x05 & (~x02 ^ x07)) | (x00 & ~x02 & ~x05 & x07))) | (x02 & ~x05 & ~x07 & x08))))) | (x01 & ~x06 & ((x08 & ((x00 & ~x07 & (x02 ? x04 : ~x05)) | (~x00 & ~x02 & ~x04 & ~x05 & x07))) | (x05 & ~x08 & ((~x00 & ~x04 & (~x07 | (x02 & x07))) | (x00 & x02 & x04 & x07))))) | (~x00 & ~x01 & x02 & x07 & ~x08 & ~x04 & ~x05))) | (~x01 & ((~x00 & ~x04 & x07 & ((~x02 & ~x05 & x06 & x08) | (x02 & x05 & ~x06 & ~x08))) | (x00 & ~x02 & x04 & ~x07 & ~x08 & x05 & x06))) | (x00 & x01 & x02 & ~x05 & x06 & (x04 ? (~x07 & x08) : (x07 & ~x08))))) | (~x03 & ((x05 & ((x06 & (x08 ? (x01 ? (((x07 ^ x10) & (x00 ? (x02 & x04) : (~x02 & ~x04))) | (~x00 & ~x02 & x04 & ~x07 & ~x10)) : ((~x00 & x02 & ~x07 & (~x04 ^ x10)) | (x00 & ~x02 & ~x04 & x07 & ~x10))) : ((x07 & ((~x02 & ((x00 & ~x10 & (~x04 | (x01 & x04))) | (~x01 & ~x04 & x10))) | (~x00 & x01 & x02 & x04 & x10))) | (~x00 & x01 & x02 & ~x07 & x10)))) | (~x06 & (x04 ? ((x07 & ((x00 & x01 & (~x08 ^ x10)) | (~x01 & x02 & ~x10 & (~x08 | (~x00 & x08))))) | (~x00 & ~x01 & ~x02 & x08 & ~x10)) : ((~x02 & ((~x00 & ~x08 & ((x07 & x10) | (x01 & ~x07 & ~x10))) | (x00 & x01 & ~x07 & x08 & x10))) | (~x00 & ~x01 & x02 & ~x07 & ~x10)))) | (~x00 & ~x01 & ~x07 & x10 & (x02 ? (x04 & ~x08) : (~x04 & x08))))) | (~x05 & (x07 ? ((x10 & (x01 ? (x06 & ((x00 & x08 & (x02 ^ x04)) | (~x02 & ~x04 & ~x08))) : (x00 ? (x06 & (x02 ? x04 : (~x04 & x08))) : (x04 & ~x06 & (x02 ^ x08))))) | (~x00 & ((x01 & ((x02 & ~x10 & (x04 ? (~x06 & x08) : x06)) | (~x02 & ~x04 & ~x06 & x08))) | (~x01 & ~x02 & x04 & x06 & x08)))) : ((x06 & ((~x01 & (x00 ? (x02 ? (~x04 & ~x08) : (x08 & x10)) : (x04 & (x02 ? ~x10 : (~x08 & x10))))) | (x00 & x01 & ~x08 & (x02 ? (~x04 & x10) : (x04 & ~x10))))) | (x00 & x01 & ~x02 & ~x04 & ~x08 & x10)))) | (x04 & ~x07 & x08 & ~x10 & ((x00 & ~x01 & x02 & x06) | (~x00 & x01 & ~x02 & ~x06))))) | (x02 & ~x04 & x00 & ~x01 & ~x05 & ~x06 & x07 & ~x08 & ~x10))) | (x09 & ((~x08 & ((~x05 & (x01 ? ((x10 & (x02 ? (x03 ? (~x06 & x07 & (~x04 | (~x00 & x04))) : ((x00 & x04 & (x06 ^ x07)) | (x06 & ~x07 & ~x00 & ~x04))) : ((x00 & x07 & (x03 ? (x04 & x06) : (~x04 & ~x06))) | (~x00 & x03 & ~x04 & ~x06 & ~x07)))) | (~x02 & x06 & x07 & ~x10 & (x00 ? (~x04 | (~x03 & x04)) : (x03 & ~x04)))) : (x00 ? ((x02 & ((x03 & ((~x04 & x06 & (x07 ^ ~x10)) | (~x07 & ~x10 & x04 & ~x06))) | (~x03 & ~x04 & ~x06 & ~x07 & x10))) | (~x02 & x03 & ~x04 & x06 & x07 & ~x10)) : (x04 ? ((~x02 & ~x03 & ~x06 & x07 & x10) | (x02 & x03 & x06 & ~x07 & ~x10)) : (x06 ? (x07 & (x02 ? ~x10 : (~x03 & x10))) : (x02 ? (x03 ? (~x07 & ~x10) : (x07 & x10)) : (x07 & (~x03 ^ x10)))))))) | (x05 & (x01 ? ((~x04 & ((~x10 & (x00 ? ((~x02 & (x03 ? (x06 & x07) : ~x07)) | (x02 & x03 & ~x06 & ~x07)) : ((x02 & x06 & (~x07 | (~x03 & x07))) | (~x02 & ~x03 & ~x06 & x07)))) | (~x03 & ~x07 & x10 & (x00 ? (x02 & ~x06) : (~x02 & x06))))) | (~x00 & x02 & x03 & x07 & x10 & x04 & x06)) : ((~x00 & (x06 ? (~x07 & ((x02 & x04 & x10) | (~x04 & ~x10 & ~x02 & x03))) : ((x07 & ((x02 & x10 & (~x03 ^ ~x04)) | (x04 & ~x10 & ~x02 & x03))) | (~x02 & ~x03 & ~x04 & ~x07 & x10)))) | (x00 & ((~x03 & ((x02 & ~x04 & x10 & (x06 ^ x07)) | (~x02 & x04 & ~x06 & x07))) | (~x02 & x03 & x04 & x06 & ~x07 & x10))) | (x06 & x07 & ~x10 & x02 & ~x03 & ~x04)))) | (x00 & ~x01 & x02 & x03 & x07 & x10 & x04 & ~x06))) | (x04 & ((x08 & (x07 ? (x02 ? ((x00 & ((x01 & ((x03 & x05 & x06) | (~x03 & ~x05 & ~x06 & ~x10))) | (~x01 & x03 & x05 & ~x06 & ~x10))) | (x05 & x06 & x10 & ~x00 & ~x01 & ~x03)) : (x01 ? ((x03 & ((x00 & (x05 ? (x06 & x10) : (~x06 & ~x10))) | (~x06 & x10 & ~x00 & ~x05))) | (x06 & ~x10 & ~x00 & x05)) : ((x00 & ((x03 & x05 & x10) | (~x03 & ~x05 & x06 & ~x10))) | (~x00 & ~x03 & x05 & ~x06 & x10)))) : ((x03 & (x00 ? (~x10 & ((x01 & ~x02 & ~x05 & x06) | (~x01 & x05 & ~x06))) : (~x06 & (x01 ? (x02 & ~x05) : (x10 & (x02 ^ ~x05)))))) | (~x00 & ~x03 & x10 & ((x01 & (x02 ? (x05 & ~x06) : (~x05 & x06))) | (~x06 & (x02 ? ~x01 : ~x05))))))) | (x00 & x01 & ~x07 & ~x10 & ((x05 & x06 & ~x02 & x03) | (~x05 & ~x06 & x02 & ~x03))))) | (x08 & ((~x04 & ((~x00 & (x03 ? ((x07 & ((x01 & ((~x02 & x06 & x10) | (x02 & ~x05 & ~x06 & ~x10))) | (~x01 & x02 & ~x05 & x06 & ~x10))) | (~x01 & x05 & ~x07 & (x02 ? (x06 & ~x10) : (~x06 ^ x10)))) : (x06 & ((~x01 & x05 & ((~x07 & x10) | (~x02 & x07 & ~x10))) | (x01 & ~x02 & ~x05 & x07 & ~x10))))) | (x00 & ((~x01 & ((~x02 & x03 & x05 & x06 & x07 & x10) | (x02 & ~x03 & ~x06 & ~x07 & ~x10))) | (x01 & ((~x03 & ((x02 & x05 & (x06 ? (x07 & x10) : (~x07 & ~x10))) | (~x02 & ~x05 & ~x06 & x07 & ~x10))) | (x06 & ~x07 & x10 & ~x02 & x03 & x05))) | (~x06 & x07 & x10 & ~x02 & x03 & ~x05))) | (~x01 & ~x02 & ~x03 & ~x05 & ~x06 & ~x07 & x10))) | (~x00 & x01 & ~x02 & x03 & ~x07 & x10 & ~x05 & x06))))) | (x02 & ~x10 & ((x01 & ((x00 & ((x03 & ~x04 & x05 & ~x06 & ~x07 & x08) | (~x03 & x04 & ~x05 & x06 & x07 & ~x08))) | (~x05 & ~x06 & ~x07 & ~x08 & ~x00 & x03 & ~x04))) | (~x00 & ~x01 & ~x03 & ~x04 & ~x05 & ~x06 & ~x07 & x08)));
  assign z01 = (~x04 & ((x09 & ((x01 & (x05 ? ((x03 & (x00 ? ((x08 & ((x02 & (x06 ? ~x10 : x07)) | (x07 & x10 & ~x02 & x06))) | (~x02 & x06 & ~x07 & ~x08 & x10)) : ((x02 & x06 & ~x07 & ~x08 & x10) | (~x02 & ~x06 & x07 & x08 & ~x10)))) | (x00 & ~x02 & ~x03 & x08 & ~x10 & x06 & ~x07)) : (x02 ? ((x07 & ((~x00 & ((x08 & x10 & ~x03 & x06) | (x03 & ~x06 & ~x10))) | (x08 & x10 & x00 & ~x03))) | (x00 & ~x07 & x10 & (x03 ? (x06 & x08) : (~x06 & ~x08)))) : (x00 ? (x03 & ((~x06 & (x07 ? (x08 & x10) : (~x08 & ~x10))) | (~x08 & ~x10 & x06 & x07))) : ((~x03 & x08 & (x06 ? (~x07 & ~x10) : (x07 & x10))) | (x03 & x06 & ~x07 & ~x08 & ~x10)))))) | (~x01 & ((~x05 & ((x02 & ((x07 & x10 & x03 & ~x06) | (~x07 & ~x10 & ~x03 & x06)) & (x00 ^ x08)) | (~x00 & ~x02 & ((~x03 & x07 & x10 & (~x08 | (x06 & x08))) | (x03 & ~x06 & ~x07 & x08 & ~x10))))) | (x05 & (x03 ? (x06 & x08 & ((~x02 & x07 & ~x10) | (x00 & ~x07 & x10))) : ((x06 & ((~x00 & x08 & (x02 ? (x07 & x10) : (~x07 & ~x10))) | (x00 & ~x02 & x07 & ~x08 & x10))) | (x00 & ~x02 & ~x06 & (x07 ? (x08 & ~x10) : (~x08 & x10)))))) | (x00 & ~x02 & ~x03 & x08 & ~x10 & ~x06 & ~x07))) | (~x00 & ~x02 & x03 & x05 & x08 & x10 & ~x06 & ~x07))) | (~x09 & ((~x03 & (x06 ? (x01 ? ((~x07 & ((~x05 & ((x00 & ~x10 & (x02 ^ ~x08)) | (x08 & x10 & ~x00 & x02))) | (~x00 & ~x02 & x05 & ~x08 & ~x10))) | (x00 & x07 & ((~x02 & x10 & (~x08 | (x05 & x08))) | (x02 & x05 & x08 & ~x10)))) : ((~x02 & ((x00 & x07 & ((x08 & x10) | (x05 & ~x08 & ~x10))) | (~x00 & ~x05 & ~x07 & ~x08 & ~x10))) | (x07 & x08 & ~x10 & ~x00 & x02 & ~x05))) : ((~x00 & (x01 ? (~x05 & ((x02 & ~x10 & (~x07 ^ x08)) | (~x02 & ~x07 & x08 & x10))) : ((~x02 & ~x05 & x07 & x08 & x10) | (x02 & x05 & ~x07 & ~x08 & ~x10)))) | (x00 & x01 & ~x02 & x05 & ~x08 & ~x10)))) | (x03 & ((x05 & ((x07 & ((x10 & (x00 ? (x02 & ((x01 & ~x06 & x08) | (x06 & ~x08))) : (x01 & ~x02 & (~x06 ^ x08)))) | (~x00 & ~x01 & ~x02 & x06 & ~x08 & ~x10))) | (~x06 & ~x07 & ~x10 & ~x00 & x01 & x02))) | (x02 & ~x05 & x08 & ((x07 & x10 & ~x01 & x06) | (~x00 & x01 & ~x06 & ~x07 & ~x10))))) | (x01 & ~x02 & x10 & ((~x00 & ~x05 & x06 & x07 & x08) | (x00 & x05 & ~x06 & ~x07 & ~x08))))) | (~x10 & ((~x05 & ~x06 & ~x07 & x08 & ~x00 & ~x01 & ~x02 & ~x03) | (x00 & x01 & x02 & x03 & x07 & ~x08 & x05 & x06))))) | (x04 & ((x09 & ((x02 & (x07 ? ((x10 & ((~x06 & ((~x08 & ((x01 & (x00 ? (~x03 ^ ~x05) : (~x03 & ~x05))) | (~x00 & ~x01 & x03 & x05))) | (~x01 & ~x03 & x05 & x08))) | (x03 & x06 & ((~x00 & x01 & x05 & x08) | (~x01 & ~x05 & ~x08))))) | (~x01 & ~x03 & x06 & ~x10 & ((~x00 & ~x05 & x08) | (x05 & ~x08)))) : ((~x06 & ((x03 & (((x01 ? (x05 & ~x08) : (~x05 & x08)) & (x00 ^ x10)) | (x00 & ~x01 & x05 & x08 & x10))) | (x00 & ~x01 & ~x03 & ~x05 & x08 & x10))) | (~x03 & x08 & ~x10 & (x00 ? (x01 & ~x05) : (~x01 & x05)))))) | (~x02 & ((x01 & (x10 ? (x00 ? (x05 & ((x06 & ~x07 & x08) | (x03 & ~x06 & ~x08))) : (x03 & ~x05 & x08 & (x06 ^ ~x07))) : (x00 ? ((~x03 & x06 & (x05 ? (x07 & x08) : ~x08)) | (x05 & ((x03 & ~x07 & x08) | (~x06 & x07 & ~x08)))) : (x03 & (x05 ? (x06 & ~x08) : (~x06 & (~x07 ^ x08))))))) | (~x00 & x10 & ((~x01 & ((x03 & ~x05 & (x06 ? (~x07 & x08) : (x07 & ~x08))) | (x05 & x06 & ~x08 & (~x07 | (~x03 & x07))))) | (~x06 & x07 & x08 & ~x03 & x05))) | (x00 & ~x01 & x03 & ~x05 & ~x08 & ~x10 & x06 & ~x07))) | (~x00 & ~x01 & x03 & x05 & ~x08 & x10 & ~x06 & ~x07))) | (~x09 & (x02 ? (x00 ? (x01 ? ((x07 & ((x03 & ~x05 & (x06 ? (~x08 & ~x10) : (x08 & x10))) | (~x03 & x05 & ~x06 & x08 & ~x10))) | (~x07 & ~x08 & ~x10 & ~x03 & x05 & x06)) : (x06 & ((~x03 & x10 & (x05 ? (~x07 & x08) : (x07 & ~x08))) | (x03 & x05 & ~x07 & ~x08 & ~x10)))) : (x01 & ((x03 & ((x05 & ((~x08 & x10 & x06 & ~x07) | (x08 & ~x10 & ~x06 & x07))) | (~x07 & x08 & x10 & ~x05 & x06))) | (~x07 & x08 & x10 & ~x03 & ~x05 & ~x06)))) : (x10 ? (x07 ? ((~x08 & (((~x01 ^ x05) & (x00 ? (~x03 & ~x06) : (x03 & x06))) | (x00 & ~x01 & x03 & x05 & ~x06))) | (~x00 & x01 & ~x03 & ~x05 & ~x06 & x08)) : ((x00 & x01 & x03 & ~x05 & (~x06 ^ x08)) | (~x00 & ~x01 & ~x03 & x05 & ~x06 & x08))) : ((~x01 & ((x05 & ~x06 & ((x00 & ~x07 & (~x03 ^ x08)) | (~x03 & x07 & x08))) | (~x00 & x03 & x06 & x07 & (~x08 | (~x05 & x08))))) | (~x00 & x01 & ~x03 & ~x07 & ~x08 & x05 & ~x06))))) | (~x00 & ~x01 & x02 & ~x03 & ~x05 & ~x06 & x07 & ~x08 & x10))) | (~x10 & (x01 ? ((~x02 & ~x06 & ((x00 & x07 & x08 & (x03 ? (~x05 & x09) : (x05 & ~x09))) | (~x00 & x03 & ~x05 & ~x07 & ~x08 & ~x09))) | (~x00 & x02 & ~x03 & x05 & x06 & x07 & x08 & x09)) : (x02 & x03 & ~x09 & ((~x00 & ~x07 & ~x08 & (x05 ^ ~x06)) | (x06 & x07 & x08 & x00 & ~x05))))) | (x00 & ~x01 & x02 & x03 & ~x05 & ~x06 & x07 & x08 & ~x09 & x10);
  assign z02 = (~x00 & ((x07 & (x08 ? ((x05 & ((~x01 & ((~x10 & ((x02 & ~x06 & (x03 ? (x04 & x09) : (~x04 & ~x09))) | (~x02 & x03 & x04 & x06 & ~x09))) | (~x02 & x04 & x06 & x10 & (~x03 | (x03 & x09))))) | (x01 & ~x09 & (x02 ? (x06 & ((~x04 & x10) | (x03 & x04 & ~x10))) : (x03 ? (x04 & x10) : (x04 ? (~x06 & ~x10) : x10)))) | (~x02 & x03 & ~x04 & x06 & x09 & x10))) | (x02 & ((x01 & ((x09 & ((x03 & ~x05 & ~x06 & (x04 ^ x10)) | (~x03 & x04 & x06 & ~x10))) | (x03 & ~x04 & ~x05 & ~x06 & ~x09 & ~x10))) | (x06 & x09 & x10 & x03 & x04 & ~x05))) | (~x02 & ~x03 & ~x05 & ~x06 & ((x01 & ((~x09 & x10) | (~x04 & x09 & ~x10))) | (~x09 & ~x10 & ~x01 & x04)))) : (x04 ? ((x09 & ((x01 & x03 & ((~x06 & x10 & ~x02 & x05) | (x02 & ~x05 & x06 & ~x10))) | (~x03 & ((~x01 & ((~x02 & ~x05 & ~x06 & x10) | (x02 & x05 & x06 & ~x10))) | (~x02 & ~x05 & ~x06 & ~x10))))) | (~x01 & ~x02 & ~x03 & ~x05 & x06 & ~x09 & ~x10)) : (x01 ? ((x03 & ((~x05 & ((x02 & (x06 ? (~x09 & ~x10) : x09)) | (~x02 & x06 & x09 & x10))) | (~x06 & ~x09 & ~x10 & ~x02 & x05))) | (x02 & ~x03 & x05 & ~x06 & x09 & x10)) : ((~x03 & ((x02 & ~x05 & (x06 ? (~x09 & x10) : (x09 & ~x10))) | (x05 & x06 & x09 & x10))) | (~x02 & x03 & x05 & x06 & ~x09)))))) | (~x07 & (x03 ? ((x09 & (x02 ? (x04 ? (~x06 & ((~x01 & (x05 ? (~x08 & x10) : (x08 & ~x10))) | (x08 & x10 & x01 & x05))) : ((~x05 & x06 & (x01 ? (~x08 ^ ~x10) : (~x08 & ~x10))) | (~x06 & ~x10 & ~x01 & x05))) : ((~x06 & ((~x08 & ((x01 & (x04 ? (~x05 & x10) : (x05 & ~x10))) | (~x01 & ~x04 & ~x05 & ~x10))) | (x05 & x08 & x10 & ~x01 & x04))) | (x05 & ~x08 & x10 & ~x01 & ~x04)))) | (~x09 & ((x02 & ((x01 & ~x06 & ((~x04 & x05 & x10) | (~x08 & ~x10 & x04 & ~x05))) | (x04 & x05 & x06 & (x08 ? ~x01 : x10)))) | (~x01 & ~x02 & ~x10 & ((~x04 & ~x05 & x06 & x08) | (x04 & x05 & ~x08))))) | (x01 & ~x02 & x04 & x05 & x06 & ~x08 & ~x10)) : (x09 ? (x02 ? ((x10 & ((x01 & x05 & x06 & (x04 ^ ~x08)) | (~x01 & x04 & ~x05 & ~x06 & ~x08))) | (~x01 & x06 & x08 & (x05 ? ~x04 : ~x10)) | (x01 & ~x04 & x05 & ~x06 & ~x08 & ~x10)) : (x10 & ((x01 & ~x08 & (x04 ? (x05 & ~x06) : (~x05 & x06))) | (~x01 & x04 & ~x05 & x06 & x08)))) : (x01 ? (x04 & ((x05 & x06 & ~x08 & ~x10) | (x02 & ~x05 & ~x06 & x08 & x10))) : (~x04 & x06 & ~x08 & (x02 ? ~x10 : (~x05 & x10))))))) | (x02 & x03 & ((~x01 & ~x04 & ~x05 & ~x08 & ~x09 & x10) | (x01 & x04 & x05 & ~x06 & x08 & x09 & ~x10))))) | (x00 & ((x10 & (x05 ? ((~x09 & (x02 ? ((~x06 & (x01 ? ((~x07 & x08 & ~x03 & ~x04) | (x07 & ~x08 & x03 & x04)) : (x07 & (x03 ? (x04 & x08) : (~x04 & ~x08))))) | (x06 & x07 & ~x08 & ~x01 & ~x03 & x04)) : (x03 ? ((x08 & ((x01 & (x04 ? (x06 & ~x07) : (~x06 & x07))) | (~x06 & ~x07 & ~x01 & x04))) | (x06 & x07 & ~x01 & x04)) : (~x07 & ((x01 & ~x06 & (x04 ^ ~x08)) | (x06 & x08 & ~x01 & ~x04)))))) | (x09 & ((~x04 & ((~x07 & ((x06 & ((x08 & (x01 ? (x02 ^ x03) : (x02 & x03))) | (~x01 & ~x02 & ~x03 & ~x08))) | (x01 & x02 & x03 & ~x06 & ~x08))) | (~x06 & x07 & x08 & ~x01 & x02 & x03))) | (x03 & x04 & ~x08 & ((~x01 & x02 & ~x06 & x07) | (x01 & ~x02 & x06 & ~x07))))) | (x01 & ~x02 & x03 & ~x07 & ~x08 & x04 & ~x06)) : ((x08 & ((~x01 & ((~x07 & ((x02 & ~x03 & x04 & x06 & x09) | (~x02 & x03 & ~x04 & ~x06 & ~x09))) | (x07 & (x02 ? (~x03 & (x06 ? x04 : x09)) : (x03 & (x04 ? ~x09 : (x06 & x09))))) | (~x02 & ~x03 & ~x04 & ~x06 & x09))) | (x07 & ((x06 & ((x01 & (x02 ? (x03 ? (~x04 & ~x09) : (x04 & x09)) : (~x04 & x09))) | (~x02 & x03 & ~x04 & ~x09))) | (x01 & x02 & ~x03 & x04 & ~x06 & ~x09))))) | (x02 & ~x08 & ((x07 & x09 & (x01 ? (x03 & x04) : (~x04 & (x03 | (~x03 & x06))))) | (~x03 & x04 & x06 & ~x07 & ~x09)))))) | (~x02 & ((~x10 & ((x01 & ((~x06 & ((~x03 & ((x04 & (x05 ? (~x07 & ~x08) : (x07 & x09))) | (~x04 & x05 & ~x07 & ~x08 & x09))) | (x03 & ~x04 & ~x05 & ~x07 & x08 & ~x09))) | (x03 & ~x04 & x06 & ((~x05 & ((x08 & x09) | (x07 & ~x08 & ~x09))) | (~x08 & x09 & x05 & ~x07))))) | (~x08 & ((~x01 & x05 & x07 & ((~x03 & ~x04 & x06 & x09) | (x03 & x04 & ~x06 & ~x09))) | (x03 & x04 & ~x05 & x06 & ~x07 & x09))) | (~x01 & ~x03 & ~x04 & x08 & (x05 ? (~x07 & ~x09) : (x06 ? x09 : (x07 & ~x09)))))) | (~x03 & x09 & ((~x06 & ~x07 & x08 & ~x01 & x04 & x05) | (x06 & x07 & ~x08 & x01 & ~x04 & ~x05))))) | (x02 & ~x10 & (x04 ? ((~x05 & ((x01 & x03 & ~x09 & ((~x07 & x08) | (x06 & x07 & ~x08))) | (~x03 & x06 & x07 & x08 & x09))) | (x01 & x03 & ~x06 & ((x05 & ~x07 & ~x08) | (x07 & x08 & ~x09)))) : ((x07 & ((x05 & ((~x03 & x06 & (x01 ? (x08 ^ x09) : (~x08 & ~x09))) | (~x01 & x03 & ~x06 & ~x08 & x09))) | (x01 & ~x05 & ~x06 & ((~x08 & ~x09) | (~x03 & x08 & x09))))) | (~x01 & ~x07 & ((x03 & x08 & ((x06 & x09) | (x05 & ~x06 & ~x09))) | (~x03 & x05 & x06 & ~x08 & x09)))))))) | (~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x08 & x09 & ~x10 & (x06 ^ ~x07));
  assign z03 = (~x07 & ((~x08 & (x04 ? ((x00 & ((((x02 & x03 & ~x05 & x10) | (~x02 & ~x03 & x05 & ~x10)) & (x01 ? (x06 & x09) : (~x06 & ~x09))) | (x01 & (x02 ? ((~x05 & ~x06 & x09 & x10) | (~x03 & x05 & x06 & ~x09 & ~x10)) : (x06 & ((x03 & x05 & x09 & x10) | (~x03 & ~x05 & ~x09 & ~x10))))) | (x06 & ((x10 & ((x02 & ((~x01 & x03 & x05) | (~x03 & ~x05 & x09))) | (~x01 & ~x02 & x09 & (x03 | (~x03 & x05))))) | (~x01 & ~x02 & x03 & x05 & ~x09 & ~x10))))) | (~x00 & ((~x05 & ((x06 & ((~x10 & ((~x01 & x02 & (~x03 ^ x09)) | (~x02 & ~x09 & (~x03 | (x01 & x03))))) | (x01 & x10 & (x02 ? (x03 & ~x09) : (~x03 & x09))))) | (x01 & ~x03 & ~x06 & x09 & ~x10))) | (~x02 & x05 & ((x01 & ~x06 & (x03 ? (~x09 & ~x10) : (x09 & x10))) | (~x01 & x03 & x06 & x09 & x10))))) | (x01 & x02 & ~x03 & x05 & ~x06 & x09 & ~x10)) : (x02 ? (x01 ? ((x00 & x09 & ((~x03 & ~x05 & ~x06 & ~x10) | (x06 & x10 & x03 & x05))) | (~x06 & ~x09 & ~x10 & ~x00 & ~x03 & x05)) : (x03 ? (x05 & ~x06 & x09 & (~x10 | (~x00 & x10))) : ((x06 & ((x00 & (x05 ? (~x09 & x10) : (x09 & ~x10))) | (~x05 & ~x09 & x10))) | (~x00 & ~x05 & ~x06 & ~x09 & ~x10)))) : ((x09 & ((x01 & ((x10 & (x00 ? (x03 ? (~x05 & ~x06) : (x05 & x06)) : (x05 & ~x06))) | (~x00 & x03 & x05 & x06 & ~x10))) | (x00 & ~x01 & ~x03 & ~x05 & x06 & x10))) | (x06 & ~x09 & x10 & ~x01 & x03 & x05))))) | (x08 & ((x04 & ((~x00 & ((~x05 & ((x01 & ((x06 & x10 & x02 & ~x03) | (~x02 & x03 & x09 & ~x10))) | (x06 & ~x09 & x10 & ~x01 & x02 & x03))) | (~x02 & ~x03 & x05 & ((~x06 & ~x09 & ~x10) | (~x01 & x09 & (~x06 ^ x10)))))) | (x09 & ((~x06 & (x01 ? ((x00 & ~x02 & (x03 ? (~x05 & x10) : ~x10)) | (x02 & x03 & x05 & x10)) : ((x05 & x10 & x02 & ~x03) | (x00 & ~x02 & x03 & ~x05 & ~x10)))) | (x00 & x03 & x05 & x06 & ~x10 & (~x01 ^ x02)))) | (x00 & x01 & ~x02 & ~x03 & x05 & x06 & ~x09 & ~x10))) | (~x04 & (x01 ? ((~x02 & ((x03 & ((x00 & x05 & x09 & (~x06 ^ x10)) | (~x00 & ~x05 & x06 & ~x09 & x10))) | (~x00 & ~x03 & x05 & ~x09 & x10))) | (x00 & x02 & x03 & x05 & x06 & ~x09 & x10)) : ((~x05 & ((~x10 & ((~x02 & (x00 ? (x03 & x06) : (~x03 & ~x06))) | (x03 & x09 & (x00 ? (~x06 | (x02 & x06)) : (x02 & ~x06))) | (~x00 & x02 & ~x03 & x06 & ~x09))) | (x00 & ~x02 & x03 & ~x06 & ~x09 & x10))) | (~x00 & x02 & x03 & x05 & x06 & ~x10)))) | (~x06 & ((~x01 & ((x00 & ~x05 & ((~x02 & ~x03 & x09 & x10) | (x02 & x03 & ~x09 & ~x10))) | (x05 & ~x09 & ~x10 & ~x00 & x02 & ~x03))) | (x00 & x01 & ~x02 & ~x03 & x05 & x09 & x10))))) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & x05 & ~x06 & x09 & ~x10))) | (x07 & ((x04 & ((x01 & (x00 ? (x03 ? ((~x09 & (x02 ? ((x05 & x06 & ~x08 & ~x10) | (~x05 & ~x06 & x10)) : (x10 & (x05 ? (x06 & ~x08) : (~x06 & x08))))) | (~x05 & x09 & x10 & (x02 ? (~x06 & x08) : ~x08))) : (~x05 & x08 & ((~x02 & x10 & (~x06 ^ ~x09)) | (x02 & x06 & x09 & ~x10)))) : ((x05 & (x02 ? (~x06 & ((x03 & x08 & x09 & x10) | (~x03 & ~x08 & ~x09 & ~x10))) : (x06 & x09 & (x03 ? (~x08 & x10) : (x08 & ~x10))))) | (x03 & ~x05 & ~x08 & ((~x02 & ~x06 & x09) | (x02 & x06 & ~x09 & ~x10)))))) | (~x01 & (x05 ? ((~x02 & ((x06 & ~x09 & ((~x00 & (x03 ? (x08 & x10) : (~x08 & ~x10))) | (x03 & x08 & ~x10))) | (x00 & ~x03 & ~x06 & x08 & x09 & x10))) | (x00 & x02 & ~x03 & ~x08 & (x09 ? x06 : ~x10))) : ((x09 & (x06 ? ((x02 & ((x00 & x10 & (~x08 | (~x03 & x08))) | (~x08 & ~x10 & ~x00 & ~x03))) | (~x00 & ~x02 & x03 & x08 & x10)) : (~x08 & ((x00 & ~x10 & (x02 ^ x03)) | (~x00 & ~x02 & x03 & x10))))) | (x03 & x06 & ~x09 & (x00 ? (~x08 & x10) : (~x10 & (x02 ^ ~x08))))))) | (x00 & x02 & x03 & x05 & x06 & x08 & ~x09 & x10))) | (~x04 & (x02 ? (x00 ? (~x09 & ((~x10 & ((x01 & ~x03 & (x05 ? (~x06 & ~x08) : (x06 & x08))) | (~x01 & x03 & x05 & ~x06 & ~x08))) | (~x01 & ~x05 & x06 & ~x08 & x10))) : ((~x08 & ((~x03 & ((~x06 & ((~x05 & (x01 ? (x09 ^ x10) : (x09 & x10))) | (~x01 & x05 & ~x09 & x10))) | (x01 & x05 & x06 & ~x09 & ~x10))) | (x03 & x05 & x06 & ~x09 & x10))) | (x01 & x08 & x10 & ((x05 & ~x06 & ~x09) | (x03 & ~x05 & x06 & x09))))) : (x00 ? ((~x08 & ((~x09 & ((~x03 & ~x05 & (x01 ? (~x06 ^ x10) : (x06 & ~x10))) | (~x01 & x03 & x05 & x06 & ~x10))) | (~x06 & x09 & x10 & ~x01 & x03 & x05))) | (x06 & x08 & ((x01 & ((x03 & ~x05 & ~x09) | (~x03 & x05 & x09 & ~x10))) | (~x01 & x03 & ~x05 & ~x09 & x10)))) : ((~x05 & ((~x09 & ((x08 & ((x01 & ~x03 & (x06 | (~x06 & x10))) | (~x06 & ~x10 & ~x01 & x03))) | (x06 & x10 & ~x01 & x03))) | (~x06 & x09 & ((x01 & x10 & (~x03 ^ x08)) | (x08 & ~x10 & ~x01 & ~x03))))) | (x01 & ~x03 & ~x06 & x08 & ~x09 & ~x10))))) | (~x05 & ~x08 & ~x10 & ((~x00 & x01 & ~x03 & (x02 ? (~x06 & ~x09) : (x06 & x09))) | (x00 & ~x01 & x02 & x03 & x06 & ~x09))))) | (~x02 & ((~x08 & ((~x09 & ((~x01 & ~x05 & ~x06 & ((x00 & ~x03 & (~x04 ^ x10)) | (~x04 & x10 & ~x00 & x03))) | (~x00 & x01 & ~x03 & x06 & ~x10 & x04 & x05))) | (x03 & ~x04 & ~x05 & x09 & ((~x01 & ~x06 & x10) | (x00 & x01 & x06 & ~x10))))) | (x00 & x03 & x08 & ~x10 & ((x01 & x04 & ~x05 & x06 & x09) | (~x01 & ~x04 & x05 & ~x06 & ~x09))))) | (x00 & x02 & ~x03 & x06 & ~x09 & ((~x01 & x04 & ~x05 & ~x08 & x10) | (x01 & ~x04 & x05 & x08 & ~x10)));
  assign z04 = (~x09 & ((~x06 & ((~x02 & (x01 ? (x05 ? ((~x03 & ((~x00 & x07 & (x04 ? (x08 & ~x10) : ~x08)) | (~x07 & ~x08 & ~x10 & x00 & x04))) | (~x00 & ~x04 & ~x07 & ~x08 & x10)) : ((x00 & ~x04 & (x03 ? (x08 & x10) : (~x08 & ~x10))) | (x04 & ~x10 & ((x03 & x07 & x08) | (~x00 & ~x07 & ~x08))))) : (x03 ? (x05 & ((x04 & ((~x08 & x10 & x00 & x07) | (x08 & ~x10 & ~x00 & ~x07))) | (x00 & ~x04 & x10 & (~x07 ^ x08)))) : (x04 ? ((x10 & ((x00 & (x05 ? (~x07 & ~x08) : (x07 & x08))) | (x07 & ~x08 & ~x00 & ~x05))) | (~x08 & ~x10 & ~x00 & x05)) : ((x07 & ~x08 & x10 & x00 & x05) | (x08 & ~x10 & ~x00 & ~x05)))))) | (x02 & ((x00 & (x03 ? ((~x05 & ((~x01 & ((~x07 & x08 & ~x10) | (x04 & x07 & ~x08 & x10))) | (x01 & x04 & ~x07 & x08 & x10))) | (~x01 & ~x04 & x05 & ~x07 & (~x08 ^ x10))) : ((x07 & ((x01 & ((x05 & x08 & ~x10) | (~x04 & ~x05 & ~x08 & x10))) | (~x01 & x04 & x05 & x08 & ~x10))) | (~x01 & x04 & ~x07 & (x05 ? (~x08 & ~x10) : (x08 & x10)))))) | (~x00 & ((x03 & (x04 ? ((x01 & x10 & (~x07 ^ x08)) | (~x07 & x08 & ~x10 & ~x01 & ~x05)) : (x01 ? (x10 & (x05 ? (~x07 & ~x08) : x08)) : (x07 & ~x10 & (x05 ^ x08))))) | (x07 & ~x08 & x10 & x01 & x04 & x05))) | (~x01 & x03 & x04 & ~x08 & x10 & x05 & ~x07))) | (x00 & x04 & ~x05 & ~x08 & ((~x07 & x10 & x01 & x03) | (x07 & ~x10 & ~x01 & ~x03))))) | (x06 & ((~x01 & ((~x04 & (x03 ? ((x00 & x02 & ~x05 & (x07 ? (x08 & x10) : ~x10)) | (~x00 & ~x02 & x05 & x08 & ~x10)) : (~x08 & (x00 ? ((x02 & x05 & (x07 ^ x10)) | (~x02 & ~x05 & ~x07 & x10)) : ((~x02 & ~x05 & x07 & x10) | (x02 & x05 & ~x07 & ~x10)))))) | (x04 & ((x00 & ((x08 & ((~x10 & ((x02 & ~x07 & (~x03 ^ ~x05)) | (~x05 & x07 & ~x02 & x03))) | (~x02 & ~x03 & x05 & x07 & x10))) | (~x03 & ~x05 & ~x07 & ~x08 & ~x10))) | (x02 & ((x07 & ((~x00 & ~x10 & (x03 ? (~x05 & x08) : (x05 & ~x08))) | (~x08 & x10 & x03 & x05))) | (~x07 & ~x08 & x10 & ~x00 & ~x03 & x05))))) | (x00 & ~x02 & x03 & ~x05 & x07 & ~x08 & x10))) | (x00 & ((x01 & (x03 ? (~x05 & ~x07 & ((~x02 & ~x10 & (x04 ^ x08)) | (x08 & x10 & x02 & ~x04))) : ((x10 & ((x02 & ((~x07 & x08 & ~x04 & x05) | (x07 & ~x08 & x04 & ~x05))) | (~x02 & x04 & x05 & ~x07 & x08))) | (x07 & x08 & ~x10 & ~x02 & x04 & x05)))) | (~x05 & x10 & ((~x02 & x03 & ~x04 & x07 & x08) | (x02 & ~x03 & x04 & ~x07 & ~x08))))) | (~x00 & x01 & ((x02 & x08 & ((x03 & (x04 ? (x07 & (x05 ^ x10)) : (x05 & ~x10))) | (~x03 & ~x04 & ~x05 & ~x07 & x10))) | (~x02 & x03 & x04 & ~x05 & x07 & ~x08 & ~x10))))) | (x00 & x03 & ~x05 & ~x07 & ~x10 & ((~x01 & ~x08 & (~x02 ^ x04)) | (x01 & x02 & x04 & x08))))) | (x09 & ((x04 & (x03 ? ((~x00 & (x10 ? (x05 ? ((~x01 & x02 & (x06 ? (x07 & ~x08) : (~x07 & x08))) | (x01 & ~x02 & x06 & ~x07 & x08)) : (~x06 & (x01 ? (x08 & (x02 ^ x07)) : (~x02 & x07)))) : ((x01 & x05 & ((~x06 & ~x08) | (~x02 & x07 & x08))) | (~x01 & x02 & x06 & ~x07 & ~x08)))) | (x00 & ((~x02 & ((~x10 & ((x08 & ((~x01 & (x05 ^ ~x06)) | (x06 & x07 & x01 & x05))) | (x01 & ~x08 & (x05 ? (x06 & ~x07) : ~x06)))) | (x01 & x07 & ~x08 & x10 & (~x06 | (x05 & x06))))) | (~x01 & x02 & x05 & x08 & ~x10 & x06 & x07))) | (x01 & ~x02 & ~x05 & ~x08 & x10 & x06 & x07)) : (x05 ? ((x08 & ((x01 & ((x02 & x10 & (x00 ? (x06 ^ ~x07) : (x06 & ~x07))) | (~x00 & ~x02 & ~x06 & ~x07 & ~x10))) | (~x06 & ~x07 & x10 & ~x00 & x02))) | (~x08 & ~x10 & x06 & x07 & ~x00 & ~x01 & ~x02)) : ((x02 & ((~x08 & ((~x00 & x01 & ~x06 & ~x07 & ~x10) | (x00 & ((~x07 & x10 & x01 & ~x06) | (x07 & ~x10 & ~x01 & x06))))) | (x07 & x08 & x10 & ~x00 & ~x01 & x06))) | (~x00 & ~x02 & x07 & x10 & (x06 ^ x08)) | (~x07 & x08 & ~x10 & x00 & ~x01 & ~x06))))) | (x03 & ((~x04 & (x00 ? ((~x08 & (x02 ? (x01 ? ((~x05 & x06 & x10) | (~x07 & ~x10 & x05 & ~x06)) : (x05 & x10 & (~x07 | (x06 & x07)))) : (~x05 & ((x06 & x07 & x10) | (~x07 & ~x10 & ~x01 & ~x06))))) | (~x01 & ~x05 & x08 & ((x07 & x10 & ~x02 & ~x06) | (~x07 & ~x10 & x02 & x06)))) : ((~x10 & (x01 ? ((~x05 & ~x06 & ~x07 & ~x08) | (x07 & x08 & ~x02 & x06)) : (x05 & x07 & x08 & (~x06 | (x02 & x06))))) | (~x08 & x10 & ~x06 & ~x07 & ~x01 & x02 & ~x05)))) | (x08 & x10 & ~x06 & ~x07 & x00 & x01 & ~x02 & x05))) | (~x04 & ((~x03 & (x05 ? (~x08 & ((x01 & ((x07 & x10 & ~x02 & ~x06) | (~x00 & x06 & (x02 ? (x07 ^ ~x10) : (~x07 & x10))))) | (~x00 & ~x01 & x02 & ~x06 & ~x07 & x10))) : ((~x02 & ((~x07 & ((~x00 & x10 & (x01 ? (~x06 & ~x08) : (x06 & x08))) | (~x08 & ~x10 & ~x01 & ~x06))) | (x07 & ~x08 & x10 & x00 & ~x01 & ~x06))) | (x00 & x02 & ((~x07 & ~x10 & ~x01 & ~x06) | (x07 & ~x08 & x10 & x01 & x06)))))) | (~x00 & x01 & x05 & x07 & ~x08 & (x02 ? (~x06 & x10) : (x06 & ~x10))))))) | (x00 & ~x02 & x03 & x04 & x05 & ~x07 & ~x10 & (x01 ? (x06 & x08) : (~x06 & ~x08)));
  assign z05 = (~x02 & ((~x08 & ((~x05 & (x00 ? (x01 ? ((x10 & ((x03 & ((x04 & x06 & ~x07 & x09) | (~x04 & ~x06 & x07 & ~x09))) | (~x03 & ~x04 & x06 & x07 & ~x09))) | (~x03 & x06 & x07 & (x04 ? (~x09 & ~x10) : x09))) : ((x10 & ((x04 & ((~x03 & x07 & (~x06 ^ x09)) | (x03 & ~x06 & ~x07 & x09))) | (x03 & ~x04 & (x06 ? (x07 & x09) : (~x07 & ~x09))))) | (~x04 & ~x07 & ~x10 & (x03 ? (~x06 & x09) : x06)))) : ((~x10 & (x01 ? ((x03 & x04 & ~x06 & x09) | (~x03 & ~x04 & x06 & ~x09)) : ((~x03 & ~x04 & (x06 ? (x07 & ~x09) : x09)) | (x03 & x04 & ~x06 & x07 & ~x09)))) | (~x01 & ((x03 & ((~x04 & ~x06 & ~x07 & (~x09 | (x09 & x10))) | (x04 & x06 & x07 & x09 & x10))) | (~x03 & ~x04 & ~x06 & ~x07 & ~x09 & x10)))))) | (x05 & ((x07 & (x04 ? ((x03 & ((x01 & ((~x00 & ~x10 & (~x06 ^ x09)) | (x00 & ~x06 & ~x09 & x10))) | (x00 & ~x01 & (x06 ? ~x09 : (x09 & x10))))) | (~x00 & ~x03 & ((~x06 & ~x09 & ~x10) | (x01 & x09 & x10)))) : (x00 ? ((x06 & x09 & x01 & x03) | (~x01 & ~x03 & ~x06 & ~x09 & ~x10)) : (x03 & x09 & x10 & (x01 ^ x06))))) | (~x06 & ((~x07 & (x03 ? (~x09 & ((x04 & x10 & ~x00 & ~x01) | (x01 & ~x04 & ~x10))) : ((~x10 & ((x00 & x04 & (~x01 ^ x09)) | (~x00 & ~x01 & ~x04 & ~x09))) | (~x09 & x10 & x01 & ~x04)))) | (x00 & ~x01 & ~x03 & x04 & x09 & x10))) | (~x00 & x01 & ~x03 & x04 & x06 & ~x07 & ~x09 & x10))) | (~x00 & ~x01 & x03 & ~x04 & x06 & ~x07 & x09 & ~x10))) | (x08 & ((~x10 & (x07 ? ((x01 & ((x03 & ((~x06 & ((~x05 & (x00 ? (~x04 ^ ~x09) : (~x04 & ~x09))) | (~x00 & ~x04 & x05 & x09))) | (x00 & x04 & x05 & x06 & x09))) | (x00 & ~x03 & ((x04 & ~x05 & ~x06 & x09) | (~x04 & x05 & x06 & ~x09))))) | (~x00 & ((~x09 & ((~x01 & x04 & ~x06 & (x03 ^ ~x05)) | (x05 & x06 & ~x03 & ~x04))) | (~x01 & x03 & ~x04 & x06 & (x05 | (~x05 & x09))))) | (x00 & ~x01 & x03 & ~x04 & x05 & ~x06 & ~x09)) : ((~x04 & ((~x03 & ((x00 & ((~x01 & ~x05 & x06 & x09) | (x01 & x05 & ~x06 & ~x09))) | (~x00 & ~x05 & ~x06 & ~x09))) | (~x00 & x03 & x09 & ((~x05 & ~x06) | (~x01 & x05 & x06))))) | (x03 & ((x04 & ((x00 & (x01 ? (x05 & ~x06) : (~x05 & ~x09))) | (~x00 & x01 & ~x06 & ~x09))) | (~x00 & ~x01 & x05 & ~x06 & x09))) | (~x00 & x01 & ~x03 & x04 & x05 & ~x06 & ~x09)))) | (x10 & ((~x06 & (x03 ? (~x07 & ((~x00 & ~x05 & (x01 ? (~x04 & x09) : ~x09)) | (x00 & x01 & ~x04 & x05 & x09))) : ((x04 & (x00 ? ((~x01 & x05 & x07 & x09) | (x01 & ~x05 & ~x07 & ~x09)) : (x01 & x09 & (~x07 | (x05 & x07))))) | (x05 & ~x07 & ~x09 & ~x00 & ~x01 & ~x04)))) | (~x01 & ((x07 & ((x03 & ((x04 & ((x00 & (x05 ? (x06 & ~x09) : x09)) | (~x00 & x05 & x06 & x09))) | (~x00 & ~x04 & ~x05 & x06 & ~x09))) | (~x05 & x06 & x09 & ~x00 & ~x03 & ~x04))) | (~x05 & x06 & ~x09 & ~x00 & ~x03 & ~x04))) | (~x00 & x01 & x03 & ~x04 & ~x05 & x06 & x07 & x09))) | (~x03 & ~x04 & ~x05 & x07 & ((~x00 & x01 & ~x06 & x09) | (x00 & ~x01 & x06 & ~x09))))) | (x00 & ~x01 & ~x03 & x04 & x05 & ~x06 & x07 & x09 & ~x10))) | (x02 & ((x06 & ((x03 & (x01 ? ((x04 & ((x00 & x05 & x07 & ~x08 & x09) | (~x00 & ~x05 & ~x07 & ~x09 & x10))) | (x00 & ~x08 & ((x05 & x07 & ~x09 & x10) | (~x04 & ~x05 & ~x07 & x09 & ~x10))) | (~x00 & ~x04 & x05 & (x07 ? (x08 & ~x10) : (~x09 & (~x10 | (x08 & x10)))))) : ((x09 & ((~x08 & ((x07 & (x00 ? (x04 ? (~x05 & ~x10) : (x05 & x10)) : (~x10 & (x04 ^ ~x05)))) | (~x05 & ~x07 & x10 & (~x00 | (x00 & x04))))) | (~x07 & x08 & ~x10 & ~x00 & x04 & ~x05))) | (x00 & ((~x04 & ((x08 & (x05 ? (~x09 & (~x10 | (x07 & x10))) : (x07 & ~x10))) | (~x05 & ~x07 & ~x08 & ~x09 & x10))) | (x08 & ~x09 & x10 & x04 & x05 & ~x07))) | (~x00 & ~x04 & x05 & x07 & ~x08 & ~x09 & ~x10)))) | (~x03 & ((x09 & ((~x08 & ((x05 & ((x01 & x04 & (x00 ? (~x07 & x10) : (x07 & ~x10))) | (~x00 & ~x01 & ((~x07 & ~x10) | (~x04 & x07 & x10))))) | (x00 & ~x04 & ~x05 & x10 & (~x01 ^ x07)))) | (x04 & x08 & ((~x01 & ((x00 & (x05 ? (~x07 & x10) : (x07 & ~x10))) | (x07 & ~x10 & ~x00 & x05))) | (~x00 & x01 & x05 & ~x07 & ~x10))))) | (x07 & ((~x09 & ((x04 & ((x00 & ((x01 & ~x05 & x08) | (~x08 & x10 & ~x01 & x05))) | (x08 & x10 & ~x00 & ~x05))) | (x05 & ~x08 & ~x10 & ~x00 & x01 & ~x04))) | (x05 & ~x08 & ~x10 & x00 & ~x01 & x04))) | (~x00 & ~x01 & ~x04 & ~x05 & x08 & ~x09 & ~x10))) | (~x00 & ~x01 & x05 & x10 & ((~x08 & x09 & ~x04 & ~x07) | (x04 & x07 & x08 & ~x09))))) | (~x06 & ((~x00 & ((x04 & (x03 ? (x01 ? (x08 & ((x07 & (x05 ? (~x09 ^ x10) : (~x09 & x10))) | (~x05 & ~x07 & x09 & x10))) : ((x08 & ~x09 & x10 & x05 & ~x07) | (~x05 & x07 & ~x08 & x09 & ~x10))) : ((~x08 & ((x01 & ~x09 & (x05 ? (x07 & ~x10) : (~x07 & x10))) | (x09 & x10 & x05 & ~x07))) | (~x05 & x08 & ((x07 & x09 & x10) | (x01 & ~x09 & ~x10)))))) | (~x04 & ((~x10 & ((~x08 & ((x01 & x07 & x09 & (~x03 ^ ~x05)) | (~x01 & x03 & x05 & ~x09))) | (~x01 & ~x03 & ~x05 & ~x07 & x08 & x09))) | (x01 & x03 & x05 & ~x07 & x09 & x10))) | (~x01 & x03 & ~x05 & ~x07 & x08 & ~x09 & ~x10))) | (x00 & (x04 ? ((x01 & ~x03 & ((x05 & ~x07 & (x08 ? x09 : (~x09 & ~x10))) | (~x05 & x07 & x08 & ~x09 & x10))) | (~x01 & x03 & ~x05 & ~x07 & x08 & x09 & x10)) : ((x10 & ((~x05 & ((~x01 & x07 & x09 & (x03 ^ x08)) | (x01 & ~x03 & ~x07 & ~x08 & ~x09))) | (x01 & x05 & ~x07 & (x03 ? (x08 & ~x09) : (~x08 & x09))))) | (~x01 & ~x05 & x07 & ~x08 & ~x10 & (x03 ^ x09))))) | (~x04 & ~x05 & x01 & x03 & ~x07 & ~x08 & x09 & ~x10))) | (~x04 & ~x05 & x08 & x09 & ((~x00 & ~x01 & x03 & ~x07 & x10) | (x00 & x01 & ~x03 & x07 & ~x10))))) | (~x09 & ((x08 & ((~x03 & ((x00 & ((~x01 & x04 & ~x05 & x06 & ~x07) | (~x06 & x07 & x10 & x01 & ~x04 & x05))) | (~x00 & ~x01 & ~x04 & x07 & ~x10 & x05 & ~x06))) | (~x00 & x01 & x03 & ~x04 & ~x05 & ~x06 & ~x07 & ~x10))) | (~x00 & x01 & x03 & ~x04 & x07 & ~x08 & ~x10 & ~x05 & x06))) | (~x00 & x01 & ~x03 & x04 & ~x05 & x06 & ~x07 & ~x08 & x09 & x10);
  assign z06 = (~x04 & ((~x00 & ((x09 & (x01 ? (x10 ? ((~x02 & x03 & x06 & ~x07 & x08) | (~x06 & x07 & ~x08 & x02 & ~x03 & x05)) : (x05 ? (x02 ? (x03 & (x06 ? (x07 ^ x08) : (x07 & x08))) : (~x03 & (x06 ? (x07 & ~x08) : (~x07 & x08)))) : ((x07 & ((x02 & x08 & (~x03 ^ x06)) | (~x06 & ~x08 & ~x02 & x03))) | (~x02 & ~x03 & x06 & ~x08)))) : (x03 ? ((~x10 & (x02 ? (x05 & ~x06 & (x07 ^ x08)) : (x06 & ((x07 & x08) | (~x05 & ~x07 & ~x08))))) | (~x07 & ~x08 & x10 & x02 & ~x05 & x06)) : ((x02 & ((x05 & x08 & x10 & (x06 ^ ~x07)) | (~x05 & ~x06 & ~x07 & ~x08 & ~x10))) | (x07 & x08 & x10 & ~x02 & ~x05 & ~x06))))) | (~x09 & ((x10 & ((x06 & ((~x08 & ((x01 & x03 & (x02 ? (x05 & ~x07) : (~x05 & x07))) | (~x01 & ~x03 & x05 & ~x07))) | (~x01 & ~x03 & x08 & (x02 ? (~x07 | (~x05 & x07)) : (x05 & ~x07))))) | (~x05 & ~x06 & ((~x01 & x02 & x07 & x08) | (x01 & ~x02 & ~x03 & ~x07 & ~x08))))) | (x02 & ~x03 & ~x10 & ((~x07 & ((~x01 & (x05 ? (~x06 & x08) : ~x08)) | (~x06 & x08 & x01 & ~x05))) | (x07 & x08 & ~x05 & x06))))) | (~x08 & x10 & ~x06 & ~x07 & ~x01 & x02 & x03 & ~x05))) | (x00 & ((x06 & (x07 ? (x05 ? ((~x02 & ((x01 & ~x03 & (x08 ? ~x09 : (x09 & x10))) | (~x08 & ~x10 & ~x01 & x03))) | (~x01 & x02 & x03 & (x08 ? (x09 & ~x10) : (~x09 & x10)))) : ((x01 & x02 & ((~x09 & x10 & ~x03 & x08) | (x03 & x09 & ~x10))) | (~x01 & ~x02 & x03 & x08 & ~x09 & ~x10))) : (x08 ? ((x03 & ((x02 & (x01 ? (x05 ? (~x09 & x10) : (x09 & ~x10)) : (x05 & ~x10))) | (~x01 & ~x02 & x05 & x09 & ~x10))) | (x01 & x02 & ~x03 & ~x05 & ~x09 & ~x10)) : ((x09 & ((~x10 & (x01 ? (x02 ? ~x05 : (x03 & x05)) : (~x05 & (x02 ^ ~x03)))) | (x02 & x10 & (x01 ? (x03 & ~x05) : (~x03 & x05))))) | (x01 & x03 & ~x09 & (x02 ? (x05 & ~x10) : (~x05 & x10))))))) | (~x06 & ((~x10 & (x01 ? ((~x07 & ((x02 & ((x03 & x05 & x08 & x09) | (~x03 & ~x05 & ~x08 & ~x09))) | (~x02 & x03 & ~x05 & x08 & ~x09))) | (~x02 & ~x03 & x07 & ~x08 & (~x09 | (x05 & x09)))) : ((~x02 & ~x03 & x07 & ((~x08 & x09) | (~x05 & x08 & ~x09))) | (x02 & x03 & ~x05 & ~x07 & x08 & x09)))) | (x02 & ((~x03 & ((x07 & ((x01 & ((x05 & ~x08 & ~x09) | (~x05 & x08 & x09 & x10))) | (~x01 & ~x05 & ~x08 & ~x09 & x10))) | (~x08 & x09 & x10 & ~x01 & ~x05 & ~x07))) | (~x01 & x03 & x05 & x07 & x08 & x09 & x10))) | (~x01 & ~x02 & ~x03 & ~x05 & x07 & ~x08 & x09 & x10))) | (~x01 & ~x02 & x03 & x05 & ~x07 & x08 & ~x09 & x10))) | (~x02 & ((~x03 & x06 & x10 & ((~x05 & ((x01 & (x07 ? (x08 & ~x09) : (~x08 & x09))) | (x08 & x09 & ~x01 & ~x07))) | (~x01 & x05 & x07 & x08 & x09))) | (~x05 & ~x06 & x01 & x03 & ~x07 & ~x08 & ~x09 & ~x10))) | (x01 & x02 & ~x03 & ~x05 & ~x06 & x07 & ~x08 & x09 & ~x10))) | (~x09 & ((x04 & ((x05 & ((x03 & (x08 ? ((~x00 & ~x01 & x02 & ~x07 & ~x10) | (x01 & ((~x00 & ((~x07 & x10 & ~x02 & x06) | (x07 & ~x10 & x02 & ~x06))) | (x00 & x02 & x06 & ~x07)))) : ((~x02 & ((~x06 & (x00 ? (x01 ? (~x07 & ~x10) : x07) : (x10 & (x01 ^ x07)))) | (x07 & x10 & x01 & x06))) | (x00 & x02 & ~x07 & (x01 ? (x06 & x10) : (~x06 & ~x10)))))) | (~x03 & (x10 ? ((x00 & ((~x01 & x02 & x06 & ~x07 & ~x08) | (x01 & x07 & x08 & (~x02 | (x02 & x06))))) | (~x01 & x02 & ~x06 & ~x07 & x08)) : ((~x07 & ((x00 & ~x08 & (x01 ? x02 : (~x02 & x06))) | (~x00 & ~x02 & ~x06 & x08))) | (~x00 & x01 & x02 & ~x06 & x07 & ~x08)))) | (x00 & x01 & ~x02 & x08 & ~x10 & ~x06 & x07))) | (~x05 & (x01 ? ((~x02 & ((x10 & ((~x07 & (x00 ^ x06) & (x03 ^ x08)) | (x07 & x08 & x03 & ~x06))) | (x07 & x08 & ~x10 & ~x00 & x03 & x06))) | (~x00 & x02 & x07 & ((~x08 & x10 & x03 & x06) | (x08 & ~x10 & ~x03 & ~x06)))) : (~x08 & ((x07 & ((x00 & x10 & (x02 ? (~x03 & x06) : (x03 & ~x06))) | (~x00 & ~x02 & ~x03 & ~x06 & ~x10))) | (x06 & ~x07 & x10 & ~x00 & x02 & x03))))) | (x00 & ~x01 & ~x02 & x03 & x08 & x10 & x06 & x07))) | (~x01 & ~x05 & x06 & x10 & ((x00 & x02 & x03 & x07 & x08) | (~x00 & ~x02 & ~x03 & ~x07 & ~x08))))) | (x09 & ((x04 & ((~x02 & ((~x10 & (x00 ? ((x08 & ((x01 & ((x03 & ~x05 & ~x06) | (x06 & ~x07 & ~x03 & x05))) | (~x01 & ~x03 & x05 & ~x06 & ~x07))) | (x06 & x07 & ~x08 & ~x01 & x03 & x05)) : ((~x01 & ~x08 & ((x03 & x07 & (x05 | (~x05 & x06))) | (x06 & ~x07 & ~x03 & ~x05))) | (x01 & ~x03 & ~x05 & x07 & x08)))) | (x10 & ((~x08 & ((x03 & ((x00 & x06 & x07 & (~x01 ^ x05)) | (~x00 & ~x01 & x05 & ~x07))) | (~x01 & ~x03 & x05 & (x07 ? ~x00 : ~x06)))) | (~x00 & ~x03 & x08 & ((x06 & x07 & x01 & x05) | (~x06 & ~x07 & ~x01 & ~x05))))) | (~x03 & ~x05 & x06 & ((x07 & x08 & ~x00 & ~x01) | (~x07 & ~x08 & x00 & x01))))) | (x02 & ((~x00 & ((x08 & ((~x03 & (x01 ? (~x05 & (x06 ? (x07 & ~x10) : x10)) : (x05 & (x06 ? (~x07 & x10) : (x07 & ~x10))))) | (x01 & x03 & x05 & ~x06 & ~x07))) | (x03 & x05 & ~x08 & ((~x07 & ~x10 & ~x01 & ~x06) | (x07 & x10 & x01 & x06))))) | (x00 & (x01 ? (~x08 & ((~x07 & x10 & ~x03 & ~x06) | (x06 & x07 & ~x10 & x03 & x05))) : (x03 & x08 & ((x06 & ~x07 & x10) | (x07 & ~x10 & x05 & ~x06))))) | (~x08 & ~x10 & x06 & ~x07 & ~x01 & ~x03 & x05))) | (~x00 & ~x01 & ((~x07 & ~x08 & x10 & ~x03 & ~x05 & ~x06) | (x03 & x05 & x06 & x07 & x08 & ~x10))))) | (~x00 & x01 & ~x02 & x03 & x05 & ~x06 & ~x07 & ~x08 & ~x10)));
  assign z07 = (x10 & ((~x03 & ((x00 & ((~x04 & ((~x06 & ((x01 & ((x08 & (x02 ? (~x05 & (~x07 | (x07 & x09))) : (~x07 & x09))) | (~x08 & ~x09 & ~x02 & x05))) | (x07 & ~x08 & ~x09 & ~x01 & x02 & x05))) | (~x05 & x06 & ((x07 & ((~x01 & x09 & (x02 ^ ~x08)) | (x02 & x08 & ~x09))) | (x01 & ~x07 & (x02 ? (~x08 & ~x09) : (x08 ^ x09))))))) | (x01 & ((x06 & ((x02 & ((~x08 & x09 & x05 & ~x07) | (x04 & ~x05 & x07 & x08 & ~x09))) | (~x07 & x08 & ~x09 & ~x02 & x04 & x05))) | (~x02 & x04 & ~x05 & ~x06 & x07 & x08 & ~x09))) | (~x01 & ((~x06 & ((~x08 & x09 & ((x02 & ((~x05 & x07) | (x04 & x05 & ~x07))) | (~x05 & ~x07 & ~x02 & x04))) | (~x02 & x08 & ~x09 & ((~x05 & ~x07) | (x04 & x05 & x07))))) | (x06 & x07 & ~x08 & ~x02 & x04 & ~x05))))) | (~x00 & (x04 ? (x01 ? ((x05 & ((x02 & ~x08 & ~x09 & (x06 ^ ~x07)) | (~x02 & x06 & ~x07 & x08 & x09))) | (~x02 & ~x05 & ~x07 & ((~x08 & x09) | (~x06 & x08 & ~x09)))) : (x07 & ((~x05 & ((x02 & x08 & (~x06 ^ ~x09)) | (~x02 & ~x06 & ~x08 & ~x09))) | (~x02 & x05 & x09 & (~x06 ^ x08))))) : ((~x02 & (x01 ? (x07 & ((x05 & x06 & ~x09) | (~x06 & x08 & x09))) : (~x07 & ((~x05 & ((~x08 & ~x09) | (x06 & x08 & x09))) | (x05 & ~x06 & ~x08 & x09))))) | (x07 & x08 & x09 & x01 & x02 & x05)))) | (~x01 & ~x02 & ~x04 & ~x05 & ~x06 & ~x07 & x08 & x09))) | (~x05 & ((x03 & ((x01 & ((x04 & ((~x06 & (x00 ? (~x07 & (x02 ? (x08 & x09) : (~x08 & ~x09))) : (x07 & (x02 ? (x08 & x09) : (x08 ^ x09))))) | (~x00 & x06 & ((~x02 & x07 & ~x08) | (x02 & ~x07 & x08 & ~x09))))) | (~x04 & ((x02 & ((x00 & ~x08 & (x06 ? (x07 & x09) : (~x07 & ~x09))) | (~x00 & x06 & ~x07 & x08 & x09))) | (~x00 & ~x02 & x06 & ~x07 & x08 & ~x09))) | (~x07 & ~x08 & x09 & ~x00 & ~x02 & ~x06))) | (~x01 & ((x07 & ((x09 & ((~x00 & ~x04 & ((~x06 & x08) | (~x02 & x06 & ~x08))) | (x00 & x02 & x04 & ~x06 & ~x08))) | (x00 & x04 & x08 & (x02 ? x06 : (~x06 & ~x09))))) | (x04 & ~x07 & ((x00 & ((~x02 & x06 & x08 & x09) | (x02 & ~x06 & ~x08 & ~x09))) | (~x00 & ~x02 & ~x06 & ~x08 & x09))))) | (~x06 & x07 & x08 & ~x09 & ~x00 & x02 & ~x04))) | (~x02 & ~x04 & ~x00 & ~x01 & x06 & x07 & x08 & ~x09))) | (x03 & x05 & ((x04 & ((~x08 & (x01 ? ((x06 & ((x00 & (x02 ? (x07 & x09) : ~x09)) | (~x00 & ~x02 & ~x07 & x09))) | (~x00 & x02 & ~x06 & x07 & ~x09)) : ((x00 & ~x02 & x06 & x09) | (~x00 & x02 & ~x06 & ~x07 & ~x09)))) | (x06 & x08 & ((x00 & ~x01 & (x02 ? (x07 & x09) : (~x07 & ~x09))) | (~x00 & x01 & x02 & x07 & x09))))) | (x01 & ((~x02 & ((x07 & (x00 ? ((~x06 & x08 & ~x09) | (~x04 & x06 & ~x08 & x09)) : (~x04 & ((~x08 & x09) | (x06 & x08 & ~x09))))) | (~x07 & ~x08 & ~x09 & ~x00 & ~x04 & ~x06))) | (x00 & x02 & ~x04 & ~x06 & ~x07 & x08 & ~x09))))))) | (~x10 & ((x02 & ((~x00 & ((x01 & ((~x05 & (x03 ? ((x08 & ((x04 & ((~x07 & x09) | (~x06 & x07 & ~x09))) | (~x04 & ~x06 & ~x07 & ~x09))) | (x04 & x06 & ~x07 & ~x08 & ~x09)) : ((~x08 & x09 & ~x04 & ~x07) | (x04 & x06 & x07 & x08 & ~x09)))) | (x03 & ~x04 & ~x06 & ((~x07 & ~x08 & ~x09) | (x05 & (x07 ? (~x08 & ~x09) : (x08 & x09))))))) | (~x01 & ((~x08 & ((x04 & ((x03 & x09 & (x05 ? (x06 & x07) : (~x06 & ~x07))) | (~x03 & ~x05 & x06 & x07 & ~x09))) | (~x03 & ~x04 & ~x07 & ~x09 & (x05 ^ ~x06)))) | (~x03 & ~x04 & x05 & ~x06 & x07 & x08 & x09))) | (~x03 & x04 & ~x05 & ~x06 & x07 & ~x08 & ~x09))) | (x00 & (x04 ? ((x01 & ((x03 & x05 & ~x06 & x07 & ~x08) | (~x05 & x06 & ~x07 & x08 & ~x09))) | (x06 & ~x08 & ((~x01 & ((x03 & (x05 ? (~x07 & ~x09) : (x07 & x09))) | (~x03 & ~x05 & ~x07 & ~x09))) | (~x03 & x05 & ~x07 & x09))) | (~x01 & x03 & ~x05 & ~x06 & ~x07 & x08 & ~x09)) : (x07 ? ((x06 & ((~x01 & ~x08 & (x03 ? (x05 & x09) : (~x05 & ~x09))) | (x01 & x03 & ~x05 & x08 & x09))) | (~x01 & ~x03 & x05 & ~x06 & ~x08)) : (x01 ? (x03 & x05 & (x06 ? (~x08 & x09) : ~x09)) : (~x03 & ~x05 & (x08 ? (~x06 ^ ~x09) : x09)))))) | (x06 & x07 & x08 & x09 & ~x01 & ~x03 & x04 & ~x05))) | (~x02 & ((~x06 & (x04 ? (x05 ? ((~x00 & x08 & x09 & (x01 ? x03 : (~x03 & x07))) | (x00 & ~x01 & ~x03 & ~x07 & ~x08 & ~x09)) : ((x03 & ((~x01 & (x00 ? (x07 ? (x08 & x09) : (~x08 & ~x09)) : (x07 ? (~x08 & ~x09) : (x08 & x09)))) | (x00 & x01 & ~x07 & x08 & ~x09))) | (x07 & ~x08 & ~x09 & x00 & x01 & ~x03))) : (x05 & ~x08 & ((x00 & ~x09 & (x03 ^ ~x07)) | (~x00 & ~x01 & ~x07 & x09))))) | (x06 & ((x04 & ((x00 & x01 & ~x03 & ~x05 & (x07 ? (x08 & x09) : (~x08 & ~x09))) | (~x00 & ~x01 & x03 & x08 & x09 & x05 & ~x07))) | (x07 & ((~x00 & ((x01 & ~x05 & ((~x03 & x08 & x09) | (x03 & ~x04 & ~x08 & ~x09))) | (~x01 & x03 & ~x04 & x05 & x08 & x09))) | (~x01 & ~x03 & x08 & x09 & (x05 ? x00 : ~x04)))))) | (~x00 & ~x01 & ~x03 & x04 & ~x05 & ~x07 & ~x08 & ~x09))) | (~x00 & ~x01 & x03 & x04 & ~x05 & ~x06 & ~x07 & x08 & ~x09))) | (~x08 & ((x01 & x05 & ((x00 & x04 & ~x06 & ~x07 & ~x09 & (x02 ^ x03)) | (~x00 & x02 & ~x03 & ~x04 & x06 & x07 & x09))) | (~x00 & ~x01 & x02 & ~x03 & x04 & ~x05 & ~x06 & x07 & x09))) | (x00 & ~x01 & ~x02 & x03 & ~x04 & ~x05 & x06 & x07 & x08 & ~x09);
  assign z08 = (x02 & ((x04 & (x08 ? (x05 ? (x09 ? ((x06 & ((x01 & ((~x00 & (x03 ? (x07 & ~x10) : (~x07 & x10))) | (~x07 & x10 & x00 & x03))) | (x00 & ~x01 & (x03 ? (x07 & ~x10) : ~x07)))) | (~x00 & ~x03 & ~x06 & (x01 ? (x07 ^ ~x10) : (~x07 & x10)))) : ((~x00 & x01 & ((x03 & ~x07 & (~x06 ^ x10)) | (x07 & ~x10 & ~x03 & x06))) | (~x06 & x07 & x10 & x00 & ~x01 & ~x03))) : (x00 ? ((x06 & ((~x01 & ((~x07 & x09 & ~x10) | (x03 & x07 & x10))) | (x01 & ~x03 & ~x07 & x09 & x10))) | (x01 & ~x06 & ((x03 & (x07 ? (x09 & x10) : (~x09 & ~x10))) | (~x03 & x07 & ~x09 & ~x10)))) : ((~x09 & ((~x07 & ((x01 & ~x03 & (~x06 ^ x10)) | (~x06 & x10 & ~x01 & x03))) | (x06 & ~x10 & ~x01 & x03))) | (~x01 & x03 & x07 & x09 & x10)))) : (x10 ? (x01 ? ((~x00 & x03 & ~x05 & x07 & x09) | (x00 & ~x03 & x05 & ~x07 & ~x09)) : ((x06 & (x00 ? ((~x03 & x05 & ~x09) | (x03 & ~x05 & x07 & x09)) : (x07 & (x03 ? x05 : (~x05 & ~x09))))) | (x00 & ~x06 & x09 & ((~x05 & ~x07) | (x03 & x05 & x07))))) : (x00 ? ((x07 & ((~x01 & x05 & ((~x06 & x09) | (x03 & x06 & ~x09))) | (~x03 & ~x05 & ((~x06 & x09) | (x01 & x06 & ~x09))))) | (x01 & ~x07 & ((x03 & ~x05 & x06 & x09) | (~x03 & (x05 ? (x06 & x09) : (~x06 & ~x09)))))) : (x05 ? ((x01 & ((x03 & x06 & ~x07 & x09) | (~x03 & ~x06 & x07 & ~x09))) | (x06 & x07 & ~x01 & ~x03)) : ((~x01 & x06 & ~x07 & (~x03 ^ x09)) | (x03 & ~x06 & x07 & ~x09))))))) | (~x04 & ((~x09 & (x10 ? ((x06 & (x03 ? ((x00 & ~x07 & (x01 ? ~x08 : (~x05 & x08))) | (~x00 & ~x01 & ~x05 & x07 & x08)) : (x00 ? (~x01 & (x05 ? (x07 ^ x08) : (~x07 & ~x08))) : (x01 & (x05 ? (x07 & x08) : ~x07))))) | (x00 & x01 & x03 & x07 & ~x08 & x05 & ~x06)) : (x00 ? (x08 & ((x01 & ((x03 & ~x07 & (x05 ^ x06)) | (~x06 & x07 & ~x03 & x05))) | (~x06 & x07 & ~x03 & ~x05))) : (x06 ? ((x01 & ~x08 & (x03 ? (~x05 & ~x07) : (x05 & x07))) | (~x01 & x03 & x05 & ~x07 & x08)) : (x01 ? (x03 & (x05 ? (~x07 & ~x08) : (x07 & x08))) : (~x03 & (x05 ? (~x07 & x08) : (x07 & ~x08)))))))) | (x09 & ((~x03 & ((x10 & (x01 ? ((~x05 & ((~x00 & ~x08 & (x06 ^ x07)) | (x07 & x08 & x00 & x06))) | (~x07 & x08 & x05 & ~x06)) : (x06 & ((x00 & x08 & (~x05 ^ x07)) | (~x07 & ~x08 & ~x00 & x05))))) | (x08 & ~x10 & ((~x00 & (x01 ? (~x06 & x07) : (~x05 & ~x07))) | (x00 & ~x01 & x05 & ~x06 & x07))))) | (~x01 & x03 & x07 & ((~x08 & (x00 ? (x05 ? x06 : (~x06 & ~x10)) : (x05 & (~x06 ^ x10)))) | (~x00 & x05 & x06 & x08 & ~x10))))) | (x00 & ~x01 & x03 & ~x05 & x08 & x10 & ~x06 & x07))) | (~x09 & ((x07 & ((x10 & ((~x00 & ((x01 & ~x03 & x05 & ~x06 & x08) | (~x01 & x03 & ~x05 & x06 & ~x08))) | (~x05 & x06 & x08 & x00 & x01 & ~x03))) | (x00 & x05 & ~x06 & ~x08 & ~x10 & (x01 ^ ~x03)))) | (x00 & x01 & x03 & x05 & x08 & x10 & x06 & ~x07))) | (~x00 & x01 & x03 & ~x05 & x06 & ~x07 & x08 & x09 & x10))) | (x00 & ((x01 & (x04 ? ((~x02 & (x03 ? ((~x08 & (((x06 ? (x07 & x09) : (~x07 & ~x09)) & (~x05 ^ x10)) | (~x05 & x06 & ~x07 & x09 & x10))) | (~x07 & x08 & x09 & (x05 ? x10 : (x06 & ~x10)))) : (x10 & ((x05 & ((~x07 & ~x08 & x09) | (x08 & (x06 ? (x07 & ~x09) : (~x07 | (x07 & x09)))))) | (~x05 & ~x06 & ~x07 & x08 & x09))))) | (x07 & ~x08 & ~x09 & ~x10 & ~x03 & x05 & ~x06)) : ((~x02 & ((x09 & ((x07 & ((~x03 & ~x06 & (x05 ? (~x08 & ~x10) : (x08 & x10))) | (x03 & ~x05 & x06 & x08 & x10))) | (x05 & x06 & ((x03 & ((~x08 & x10) | (~x07 & x08 & ~x10))) | (~x08 & ~x10 & ~x03 & ~x07))))) | (x03 & x08 & ~x09 & ((~x06 & ~x07 & x10) | (~x05 & x07 & (~x06 ^ ~x10)))))) | (~x08 & ~x09 & ~x10 & ~x05 & ~x06 & x07)))) | (~x01 & ((~x10 & ((~x02 & ((x09 & ((x06 & ((x07 & (x03 ? (~x08 & (x04 ^ ~x05)) : (x04 & ~x05))) | (~x03 & ~x04 & ~x05 & ~x07 & ~x08))) | (~x04 & ~x05 & ~x06 & (x03 ? (~x07 ^ x08) : (~x07 & x08))))) | (~x06 & ~x07 & ~x08 & ~x09 & (x03 ? ~x05 : (~x04 & x05))))) | (x03 & x04 & ((~x05 & x06 & x07 & x08 & x09) | (x05 & ~x06 & ~x07 & ~x08 & ~x09))))) | (~x02 & x10 & ((x06 & ((~x03 & ((x04 & ((x05 & x08 & x09) | (~x05 & x07 & ~x08 & ~x09))) | (~x04 & x05 & ~x07 & ~x08 & ~x09))) | (x03 & ~x04 & x05 & x07 & x08 & x09))) | (x03 & x04 & ~x05 & ~x09 & ((~x06 & x07 & x08) | (~x07 & ~x08))))))) | (~x02 & ~x04 & ~x05 & x06 & ~x10 & ((~x03 & x07 & x08 & x09) | (~x08 & ~x09 & x03 & ~x07))))) | (~x02 & ((~x00 & ((x07 & ((~x04 & (x01 ? ((x09 & (x08 ? ((x06 & (x03 ? (~x05 ^ x10) : x10)) | (~x06 & ~x10 & ~x03 & x05)) : (x10 & (x05 ? x03 : x06)))) | (~x03 & ~x05 & x08 & ~x09 & ~x10)) : ((~x10 & ((x03 & ~x09 & (x05 ? (x06 & ~x08) : (~x06 & x08))) | (~x03 & ~x05 & ~x06 & ~x08 & x09))) | (~x03 & x09 & x10 & (x05 ? (~x08 | (x06 & x08)) : (~x06 & x08)))))) | (x04 & ((x09 & ((~x06 & ((~x01 & ~x10 & (x03 ? (x05 & ~x08) : (~x05 & x08))) | (~x05 & x08 & x10 & x01 & ~x03))) | (x01 & ~x03 & x06 & x10 & (~x05 ^ x08)))) | (x01 & ~x09 & ((~x03 & x06 & (x05 ? (~x08 & x10) : (x08 & ~x10))) | (x03 & ~x05 & ~x06 & x08 & ~x10))))) | (x01 & x03 & x05 & x06 & x08 & ~x09 & ~x10))) | (~x07 & (x03 ? (x08 & ((x05 & ((x01 & (x04 ? (x06 ? (x09 & ~x10) : (~x09 & x10)) : (~x06 & ~x10))) | (~x06 & x09 & ~x10 & ~x01 & ~x04))) | (x04 & ~x05 & ~x09 & ~x10))) : ((x06 & ((~x08 & ((x01 & ((~x04 & x05 & ~x09 & x10) | (x04 & ~x05 & x09 & ~x10))) | (~x01 & x04 & ~x05 & x09 & x10))) | (~x01 & x04 & x08 & ~x10 & (x05 ^ x09)))) | (~x04 & x08 & ((x01 & ((~x06 & ~x09 & ~x10) | (~x05 & x09 & x10))) | (~x01 & ~x05 & ~x06 & ~x09 & x10)))))) | (~x04 & ~x05 & x01 & x03 & ~x06 & ~x08 & x09 & x10))) | (~x01 & ~x04 & x06 & x08 & ~x09 & ((~x07 & x10 & x03 & x05) | (x07 & ~x10 & ~x03 & ~x05))) | (x01 & ~x03 & x04 & x05 & ~x06 & ~x07 & ~x08 & x09 & ~x10))) | (~x00 & ~x04 & x05 & ~x06 & ~x07 & ~x09 & x10 & (x01 ? (~x03 & ~x08) : (x03 & x08)));
  assign z09 = (x08 & ((x07 & ((~x05 & (x04 ? (x00 ? ((x09 & ((x01 & x03 & (x02 ? (~x06 & x10) : (x06 & ~x10))) | (~x01 & ~x02 & ~x03 & ~x06 & x10))) | (~x01 & ~x03 & ~x09 & ((x06 & ~x10) | (x02 & ~x06 & x10)))) : ((~x03 & ((~x02 & ((x06 & ~x09 & x10) | (x09 & ~x10 & ~x01 & ~x06))) | (x01 & x02 & x06 & x10))) | (~x01 & x02 & x03 & ~x10 & (~x06 ^ ~x09)))) : ((~x06 & (x00 ? ((~x01 & ((~x02 & ~x03 & (x09 ^ x10)) | (x02 & x03 & x09 & x10))) | (x01 & ~x02 & ~x03 & ~x09 & ~x10)) : (x01 ? (~x10 & (x02 ? (~x03 & ~x09) : (x03 & x09))) : (x02 & (x03 ? (~x09 & x10) : x09))))) | (~x00 & ~x01 & ~x02 & ~x03 & x06 & x09 & ~x10)))) | (x05 & ((x03 & ((~x01 & (x00 ? (x10 & ((x02 & (x04 ? (~x06 & ~x09) : (x06 & x09))) | (~x02 & ~x04 & ~x06 & ~x09))) : (~x10 & ((~x02 & x09 & (~x06 | (~x04 & x06))) | (x02 & ~x04 & x06 & ~x09))))) | (~x00 & ((x04 & ~x09 & ((~x02 & x06 & x10) | (x01 & x02 & ~x06 & ~x10))) | (x01 & x02 & x09 & ((x06 & ~x10) | (~x04 & ~x06 & x10))))))) | (~x00 & ~x03 & (x06 ? (x09 & ((x02 & ~x04 & x10) | (~x01 & ~x02 & x04))) : (~x09 & ((x01 & x10 & (~x02 ^ x04)) | (~x01 & x02 & x04 & ~x10))))))) | (~x00 & x01 & ~x02 & ~x03 & ~x04 & x06 & ~x09 & ~x10))) | (x00 & ((~x01 & ((x03 & ((~x06 & ~x10 & ((x02 & ~x09 & (x04 ? (x05 & ~x07) : ~x05)) | (~x02 & ~x04 & x05 & ~x07 & x09))) | (x05 & x06 & ~x07 & x10 & (x09 ? ~x04 : ~x02)))) | (~x02 & ~x03 & x06 & ~x07 & ((~x04 & x05 & ~x09) | (x04 & ~x05 & x09 & x10))))) | (~x07 & ((x01 & (x02 ? ((x03 & ~x05 & ((~x04 & ~x06 & x09 & x10) | (x04 & x06 & ~x09 & ~x10))) | (x05 & ((~x04 & x06 & x09 & x10) | (~x03 & ~x06 & ~x09 & ~x10)))) : ((~x03 & ((~x04 & x05 & ~x06 & x09 & ~x10) | (x04 & ~x05 & x06 & ~x09 & x10))) | (~x06 & x09 & ~x10 & x03 & x04 & x05)))) | (x05 & x06 & x09 & x10 & x02 & ~x03 & x04))))) | (~x07 & ((~x00 & (x01 ? (x02 ? (x03 & ~x06 & (x04 ? (x09 & x10) : (x05 ? (~x09 & x10) : (x09 & ~x10)))) : ((~x09 & ((~x03 & x04 & x06 & ~x10) | (~x05 & ~x06 & (x03 ? (x04 ^ x10) : (~x04 & ~x10))))) | (x03 & x04 & x06 & x09 & ~x10))) : ((x06 & ((x04 & x10 & ((x02 & x05 & (~x03 ^ x09)) | (~x02 & x03 & ~x05 & x09))) | (x02 & ~x03 & ~x04 & ~x05 & ~x09 & ~x10))) | (x05 & ~x06 & ((~x02 & x10 & ((~x04 & x09) | (~x03 & x04 & ~x09))) | (x02 & x03 & ~x04 & x09 & ~x10)))))) | (x02 & x05 & ((x01 & x06 & x09 & ~x10 & (~x03 ^ ~x04)) | (~x01 & ~x03 & ~x04 & ~x09 & x10))))) | (~x00 & x01 & x02 & x03 & ~x04 & ~x05 & ~x06 & ~x09 & ~x10))) | (~x08 & ((~x06 & (x04 ? (x09 ? ((x00 & ((x05 & ((x10 & ((x01 & (x02 ? (x03 & ~x07) : x07)) | (~x01 & ~x02 & x03 & x07))) | (~x01 & x02 & x03 & ~x10))) | (x01 & ~x02 & ~x03 & ~x07 & (~x10 | (~x05 & x10))))) | (~x02 & x03 & ~x05 & ~x10 & ((x01 & x07) | (~x00 & ~x01 & ~x07)))) : ((x02 & (x00 ? ((~x07 & x10 & x01 & x03) | (~x01 & ~x03 & ~x05 & ~x10)) : (x05 & x10 & (x01 ? (x03 ^ ~x07) : (~x03 & x07))))) | (~x01 & ((~x02 & ((~x03 & ((~x05 & x07 & ~x10) | (x00 & x10 & (x05 ^ x07)))) | (~x00 & x03 & x05 & x07 & ~x10))) | (~x00 & x03 & ~x05 & x07 & x10))) | (~x00 & x01 & ~x10 & ((~x03 & ~x05 & x07) | (~x02 & x03 & x05 & ~x07))))) : (x02 ? ((~x01 & ((~x07 & ((x00 & x10 & (x03 ? (x05 & ~x09) : x09)) | (x03 & x05 & ~x09 & ~x10))) | (~x00 & ~x05 & x07 & x09 & x10))) | (~x00 & ((x01 & x07 & ((~x03 & x05 & ~x09 & x10) | (x03 & ~x05 & x09 & ~x10))) | (~x07 & ~x10 & ~x03 & x05))) | (x01 & ~x03 & x05 & x07 & ~x10)) : ((x03 & ((x07 & ((~x00 & ~x10 & (x01 ? (x05 & x09) : (~x05 & ~x09))) | (x00 & ~x01 & ~x05 & x09 & x10))) | (x00 & ~x07 & (x01 ? (x09 & (~x05 ^ x10)) : (~x05 & ~x09))))) | (x00 & x01 & ~x05 & ~x07 & ~x09 & ~x10))))) | (x06 & ((x00 & (x07 ? ((x02 & (x01 ? (x03 & ((~x04 & ~x05 & x09 & x10) | (x04 & x05 & ~x10))) : (x09 & ((x04 & ~x05 & ~x10) | (~x03 & ~x04 & x05 & x10))))) | (~x01 & x03 & ~x04 & x10 & ((~x05 & ~x09) | (~x02 & x05 & x09)))) : (x01 ? ((~x05 & ((x02 & ~x04 & (x03 ? (~x09 & x10) : (x09 & ~x10))) | (~x02 & x03 & x04 & x09 & ~x10))) | (x05 & ~x09 & x10 & ~x02 & ~x03 & x04)) : ((x02 & ((x03 & ~x04 & ~x10 & (x05 ^ ~x09)) | (~x03 & x04 & x05 & ~x09 & x10))) | (~x03 & ~x04 & ~x05 & ~x09 & ~x10))))) | (~x00 & (x05 ? ((x02 & ((x03 & ((x01 & x09 & x10 & (x04 ^ x07)) | (~x01 & ~x04 & ~x07 & ~x09 & ~x10))) | (~x01 & ~x03 & x04 & x07 & x09 & ~x10))) | (~x09 & ((x01 & ((~x04 & ((x03 & x07 & ~x10) | (~x02 & x10 & (x03 ^ x07)))) | (~x02 & ~x03 & x04 & x07 & ~x10))) | (~x01 & ~x02 & ~x03 & ~x04 & x07)))) : ((x09 & ((~x04 & ((x07 & ((x01 & ~x02 & (~x10 | (~x03 & x10))) | (~x01 & x02 & x03 & x10))) | (~x01 & x02 & ~x03 & ~x07 & x10))) | (~x01 & x02 & ~x03 & x04 & ~x10))) | (~x01 & x02 & x03 & x04 & x07 & ~x09 & x10)))) | (~x01 & ~x02 & x03 & x04 & ~x05 & x07 & x09 & ~x10))) | (~x10 & ((x00 & x02 & x04 & ((x01 & ~x03 & x05 & ~x07 & x09) | (~x01 & x03 & ~x05 & x07 & ~x09))) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ~x07 & ~x09))))) | (~x05 & ((~x00 & x10 & ((~x01 & ~x03 & x04 & x09 & (x02 ? (x06 & x07) : (~x06 & ~x07))) | (~x04 & ~x06 & x07 & ~x09 & x01 & x02 & x03))) | (x00 & ~x01 & ~x02 & x03 & x04 & x06 & ~x07 & ~x09 & ~x10)));
  assign z10 = (x08 & ((x04 & ((~x00 & (x03 ? ((x07 & ((x05 & ((~x01 & ((x06 & ~x09 & ~x10) | (~x02 & x10 & (~x06 ^ x09)))) | (~x02 & ~x06 & x09 & (~x10 | (x01 & x10))))) | (x02 & ~x05 & x10 & (x01 ? (~x06 ^ x09) : (x06 & ~x09))))) | (~x05 & ~x07 & ((x06 & ((~x01 & (x02 ? (x09 & ~x10) : x10)) | (x01 & ~x02 & ~x09 & ~x10))) | (~x02 & ~x06 & x09 & ~x10)))) : ((~x07 & ((~x01 & ((~x05 & x06 & ~x09 & x10) | (x09 & ~x10 & ~x02 & x05))) | (~x06 & x09 & ~x10 & x01 & x02 & x05))) | (x01 & ~x02 & ((~x05 & ~x06 & ~x09 & x10) | (x05 & x06 & x07 & x09 & ~x10)))))) | (x00 & (x07 ? (x01 ? (x02 ? (~x03 & (x05 ? (x06 & x09) : (~x09 & ~x10))) : (x03 & x05 & (x06 ? (x09 & ~x10) : x10))) : ((x09 & (x02 ? ((~x05 & ~x06 & (~x10 | (x03 & x10))) | (~x03 & x05 & ~x10)) : ((~x03 & ~x05 & x06) | (~x06 & x10 & x03 & x05)))) | (~x05 & ~x09 & x10 & (x02 ? (~x03 & ~x06) : (x03 & x06))))) : ((x06 & (x01 ? (x05 & ((~x02 & x10 & (~x03 ^ x09)) | (x02 & ~x03 & ~x09 & ~x10))) : ((x10 & ((x02 & x09 & (x03 ^ ~x05)) | (~x02 & x03 & x05 & ~x09))) | (x02 & ~x03 & ~x05 & ~x09 & ~x10)))) | (~x02 & x03 & ~x05 & ~x06 & ~x09 & x10)))) | (~x01 & x02 & x03 & x05 & x06 & x07 & x09 & ~x10))) | (~x04 & ((x03 & (x02 ? ((~x06 & ((x10 & (x00 ? (~x05 & (x01 ? (x07 & x09) : (~x07 & ~x09))) : (x05 & x07 & (x01 | (~x01 & x09))))) | (~x07 & x09 & ~x10 & x00 & x01 & x05))) | (x00 & ~x05 & x06 & ((~x01 & (x07 ? (~x09 & x10) : (x09 & ~x10))) | (x09 & ~x10 & x01 & x07)))) : (x00 ? ((~x01 & ((x05 & ~x07 & x10 & (~x06 ^ x09)) | (~x05 & x06 & x07 & x09 & ~x10))) | (x06 & ~x07 & x10 & x01 & ~x05)) : ((x10 & (x01 ? (x06 & (x05 ? (~x07 & x09) : (x07 & ~x09))) : (~x06 & x09 & (x05 | (~x05 & x07))))) | (x05 & ~x10 & ((~x01 & x06 & ~x07 & x09) | (x07 & ~x09 & x01 & ~x06))))))) | (~x03 & (x05 ? ((x00 & ((~x01 & ~x09 & ((~x02 & x07 & x10) | (~x07 & ~x10 & x02 & ~x06))) | (~x07 & x09 & ~x10 & x01 & x02 & x06))) | (~x00 & ((x01 & ((~x07 & ~x10 & x02 & x06) | (~x02 & x07 & ~x09 & x10))) | (x07 & x09 & x10 & ~x01 & x02 & x06))) | (x07 & x09 & ~x10 & x01 & ~x02 & x06)) : ((x09 & ((~x02 & ((~x00 & ((x01 & (x06 ? (x07 & x10) : (~x07 & ~x10))) | (x07 & ~x10 & ~x01 & ~x06))) | (x00 & ~x01 & x06 & ~x07 & x10))) | (x00 & x02 & ((x06 & x07 & ~x10) | (~x07 & x10 & x01 & ~x06))))) | (~x00 & ~x01 & ~x02 & ~x06 & ~x07 & ~x09 & ~x10)))) | (x00 & ~x01 & x02 & ~x05 & x07 & ~x09 & ~x10))) | (~x00 & x05 & x06 & ~x07 & ~x10 & ((x01 & ~x02 & ~x03 & x09) | (~x01 & x02 & x03 & ~x09))))) | (~x08 & (x10 ? ((x06 & (x00 ? (x03 ? ((x02 & ((x01 & x05 & (x04 ? (x07 & x09) : (~x07 & ~x09))) | (~x01 & ~x05 & x07 & ~x09))) | (~x01 & ~x02 & ((x05 & ~x07 & x09) | (x04 & x07 & ~x09)))) : ((x01 & ((x02 & ~x04 & ((x07 & ~x09) | (x05 & ~x07 & x09))) | (x04 & x05 & ~x07 & ~x09))) | (~x01 & ~x04 & ~x05 & ~x07 & x09))) : ((x02 & ((~x04 & ((~x03 & ((x01 & ~x05 & (x07 ^ ~x09)) | (~x01 & x05 & ~x07 & ~x09))) | (~x01 & x03 & x05 & ~x07 & x09))) | (x03 & x04 & x05 & ~x07 & ~x09))) | (x01 & ~x02 & ~x03 & ((~x04 & ~x05 & ~x07 & x09) | (x04 & x05 & x07 & ~x09)))))) | (~x06 & ((~x04 & ((~x03 & x05 & (x00 ? (~x02 & (x01 ? (x07 & ~x09) : (~x07 & x09))) : (x02 & ~x09 & (x01 ^ x07)))) | (x01 & ~x05 & ((x00 & x02 & ~x07 & x09) | (~x02 & x03 & x07 & ~x09))))) | (~x00 & ((x03 & ((x01 & ~x09 & (x02 ? (x05 & x07) : (x04 & ~x05))) | (~x05 & x07 & x09 & ~x01 & x02 & x04))) | (~x01 & ~x02 & ~x03 & x04 & x05 & x07 & x09))) | (x04 & x05 & x07 & x09 & x00 & ~x01 & x02 & ~x03))) | (~x00 & x01 & ~x02 & x03 & x04 & ~x05 & ~x07 & x09)) : ((x09 & ((x00 & (x06 ? (~x07 & ((x02 & ((x01 & ((x03 & ~x04 & ~x05) | (x04 & x05))) | (~x01 & x03 & x04 & x05))) | (~x01 & ~x02 & x03 & x04 & ~x05))) : (x02 ? (x03 & ((x01 & x04 & (~x05 ^ x07)) | (~x05 & ~x07 & ~x01 & ~x04))) : (x01 ? (~x03 & ~x04) : (x07 & (x03 ? (~x04 & ~x05) : (x04 & x05))))))) | (~x00 & ((~x06 & ((x01 & x07 & ((~x02 & ~x03 & ~x04 & x05) | (x02 & x03 & x04 & ~x05))) | (~x02 & ~x03 & x04 & ~x05) | (~x01 & x02 & x03 & ~x04 & x05 & ~x07))) | (~x01 & x03 & ~x05 & x06 & x07 & (x02 ^ x04)))) | (~x01 & ~x02 & ~x03 & x06 & ~x07 & x04 & x05))) | (~x09 & ((~x01 & (x05 ? ((~x07 & ((~x00 & ((x04 & x06 & x02 & ~x03) | (~x04 & ~x06 & ~x02 & x03))) | (x00 & x02 & x03 & ~x04 & x06))) | (x00 & ~x02 & ((x03 & x04 & x06) | (~x03 & ~x04 & ~x06 & x07)))) : ((x02 & ((x00 & ((x03 & x04 & x07) | (~x04 & x06 & ~x07))) | (~x00 & x03 & x04 & x06 & x07))) | (~x04 & ~x06 & ~x07 & x00 & x03)))) | (x00 & x01 & ((x05 & ((x02 & x06 & (x03 ? (x04 & x07) : ~x04)) | (~x02 & ~x03 & ~x06 & ~x07))) | (~x05 & x06 & ~x07 & ~x02 & ~x03 & ~x04))))) | (~x00 & ~x01 & ~x02 & x03 & ~x06 & ~x07 & x04 & ~x05)))) | (~x00 & x02 & x04 & ~x10 & ((x06 & ~x07 & x09 & ~x01 & ~x03 & ~x05) | (~x06 & x07 & ~x09 & x01 & x03 & x05)));
  assign z11 = (x04 & ((~x00 & ((x02 & ((x06 & (x03 ? ((x08 & ~x09 & x10 & x05 & ~x07) | (~x05 & ((~x08 & x10 & x01 & ~x07) | (x08 & ~x09 & ~x10 & ~x01 & x07)))) : ((~x10 & ((~x05 & (x01 ? (x07 & (x08 ^ x09)) : (~x08 & x09))) | (~x01 & x05 & x07 & ~x08 & x09))) | (x08 & ~x09 & x10 & x01 & x05 & x07)))) | (~x06 & ((~x10 & (x01 ? ((x03 & x05 & ~x07 & x08 & x09) | (~x03 & ~x05 & x07 & ~x08 & ~x09)) : (~x05 & ~x08 & x09 & (x03 ^ x07)))) | (~x01 & x05 & x08 & x10 & (x03 ? (~x07 & x09) : (x07 & ~x09))))) | (~x01 & x03 & x05 & ~x07 & x08 & ~x09 & ~x10))) | (~x02 & (x01 ? (x07 & ((~x03 & ((~x05 & x09 & ((~x08 & x10) | (~x06 & x08 & ~x10))) | (x08 & x10 & x05 & ~x06))) | (x03 & ~x05 & ~x08 & ~x09 & x10))) : (x03 ? ((~x10 & ((~x05 & ~x06 & ~x07 & x08 & x09) | (x07 & ((x05 & (x06 ? x08 : (~x08 & ~x09))) | (~x05 & x06 & ~x08 & ~x09))))) | (~x05 & ~x07 & x10 & (x06 ? ~x09 : (~x08 & x09)))) : ((~x06 & ((x10 & ((x07 & ~x08 & ~x09) | (x05 & x09 & (x07 ^ x08)))) | (~x05 & x07 & x08 & ~x09 & ~x10))) | (~x05 & ~x07 & ~x08 & ~x09 & ~x10))))) | (~x01 & x05 & x06 & ~x07 & ~x10 & (x03 ? (~x08 & x09) : (x08 & ~x09))))) | (x00 & (x06 ? (x03 ? ((~x05 & ((~x08 & ((x07 & ((x01 & (x02 ? (x09 & x10) : (~x09 & ~x10))) | (~x01 & ~x02 & ~x09 & x10))) | (~x01 & x02 & ~x07 & ~x10))) | (x01 & x08 & ((~x02 & (x07 ? (x09 & ~x10) : (~x09 & x10))) | (x02 & x07 & ~x09 & ~x10))))) | (~x08 & x09 & x10 & x01 & x02 & ~x07)) : (x02 ? ((~x01 & ~x05 & ~x08 & ~x09 & x10) | (x08 & ((x05 & ((x01 & (x07 ? (~x09 & ~x10) : (x09 & x10))) | (x09 & x10 & ~x01 & x07))) | (~x01 & ((~x07 & ~x09 & ~x10) | (~x05 & x07 & x10)))))) : ((~x08 & (x01 ? (x05 & (x07 ? x10 : (~x09 & ~x10))) : (~x05 & x07 & (~x09 ^ x10)))) | (~x07 & x09 & ~x10 & (x05 ? ~x01 : x08))))) : (x10 ? ((~x02 & ((x03 & (x01 ? (x05 & (x07 ? (~x08 & x09) : (x08 & ~x09))) : (~x05 & (x07 ? (x08 & x09) : (~x08 & ~x09))))) | (x01 & ~x03 & ~x05 & x08 & (x07 ^ ~x09)))) | (~x09 & ((x01 & ((~x05 & x08 & x02 & x03) | (~x07 & ~x08 & ~x03 & x05))) | (x02 & ~x03 & ~x05 & x07 & ~x08))) | (x07 & x08 & x09 & ~x01 & x02 & x05)) : (x02 ? (x08 & ((~x01 & ~x05 & (x03 ? ~x09 : (x07 & x09))) | (x03 & x05 & x07 & x09))) : (~x03 & x05 & x07 & ~x08 & (~x09 | (x01 & x09))))))) | (~x06 & x07 & ~x08 & x09 & ~x10 & ~x01 & ~x02 & ~x03 & x05))) | (~x04 & ((x08 & ((~x02 & (x05 ? ((~x01 & ((~x03 & ((~x00 & ((~x06 & ~x07 & ~x09 & ~x10) | (x06 & x07 & x09 & x10))) | (~x09 & x10 & x00 & x07))) | (x00 & x03 & ~x10 & (x06 ? (~x07 & ~x09) : (x07 & x09))))) | (x00 & ((x01 & x07 & ~x09 & ((x06 & ~x10) | (x03 & ~x06 & x10))) | (x03 & ~x06 & ~x07 & x09 & x10))) | (~x00 & x01 & ~x03 & ~x06 & x07 & x09 & x10)) : ((~x03 & ((x07 & ((~x00 & ((~x06 & ~x09 & x10) | (x09 & ~x10 & x01 & x06))) | (x00 & ~x01 & x06 & x09 & x10))) | (x00 & ~x07 & (x01 ? (~x06 & ~x09) : (x06 & ~x10))))) | (x03 & ((x07 & ((x00 & ((~x01 & x06 & ~x10) | (x09 & x10 & x01 & ~x06))) | (~x00 & x01 & ~x06 & x09 & ~x10))) | (~x00 & ~x01 & x06 & ~x07 & x09 & x10))) | (x00 & ~x01 & ~x06 & ~x07 & x09 & ~x10)))) | (x02 & (x00 ? ((~x07 & ((~x06 & ((x01 & ~x09 & ((x05 & ~x10) | (~x03 & ~x05 & x10))) | (~x01 & x03 & ~x05 & x09 & x10))) | (~x01 & x05 & x06 & x09 & ~x10))) | (x01 & x07 & ((~x10 & ((x03 & x05 & (~x06 ^ x09)) | (~x05 & ~x06 & x09))) | (~x03 & ~x05 & x06 & ~x09 & x10)))) : ((x07 & ((x05 & (x01 ? ((x03 & x06 & ~x09) | (~x03 & ~x06 & x09 & ~x10)) : (x06 & (x03 ? (x09 & ~x10) : (~x09 & x10))))) | (~x01 & ~x05 & x10 & (x03 ? (~x06 & ~x09) : (x06 & x09))))) | (~x01 & ~x05 & x06 & ~x10 & (x03 ? ~x07 : x09))))) | (~x00 & x01 & ~x03 & ~x05 & ~x06 & x07 & x09 & ~x10))) | (~x08 & (x00 ? ((~x01 & ((x09 & (x02 ? (x07 & ((~x03 & ~x05 & ~x06 & ~x10) | (x06 & x10 & x03 & x05))) : (~x07 & ~x10 & (x03 ? (x05 & ~x06) : x06)))) | (~x06 & ((~x07 & (x02 ? ((x03 & ~x05 & x10) | (~x03 & x05 & ~x09 & ~x10)) : (~x05 & ~x09 & (x03 ^ x10)))) | (~x02 & x03 & x05 & x07 & ~x09))))) | (x06 & ((x09 & ((x01 & (x02 ? (x07 & (x03 ? (~x05 & ~x10) : x10)) : (x03 & ~x07 & (x05 ^ x10)))) | (~x02 & ~x03 & x10 & (~x05 ^ x07)))) | (~x05 & x07 & ~x09 & ~x10 & x01 & ~x02 & ~x03))) | (x01 & x02 & x03 & ~x05 & ~x06 & ((~x09 & ~x10) | (~x07 & x09 & x10)))) : ((x01 & ((x09 & ((~x06 & x07 & x10 & ~x02 & x03 & ~x05) | (x06 & ((x02 & ((~x07 & x10 & ~x03 & ~x05) | (x07 & ~x10 & x03 & x05))) | (~x02 & ~x03 & x05 & x07 & ~x10))))) | (~x03 & ~x09 & ((x02 & ~x07 & ((x06 & ~x10) | (x05 & ~x06 & x10))) | (x06 & x10 & ~x02 & x05))))) | (~x01 & ((~x03 & ((~x07 & ((x02 & ~x06 & (x09 ? ~x05 : ~x10)) | (x06 & x09 & x10 & ~x02 & x05))) | (x07 & ~x09 & x10 & ~x02 & x05 & x06))) | (x02 & x03 & ~x05 & ~x06 & x07 & ~x09 & ~x10))) | (x06 & x07 & x09 & x10 & ~x02 & ~x03 & ~x05)))) | (~x00 & x01 & ~x02 & x03 & x05 & ~x06 & ~x07 & x09 & x10))) | (x01 & x05 & ~x07 & ((~x08 & ((x00 & x06 & ~x09 & (x02 ? (~x03 & ~x10) : (x03 & x10))) | (~x06 & x09 & ~x10 & ~x00 & x02 & ~x03))) | (~x00 & x02 & x03 & ~x06 & x08 & ~x09 & ~x10))) | (~x06 & x07 & x08 & ~x09 & x10 & x00 & ~x01 & ~x02 & x03 & ~x05);
  assign z12 = (x08 & (x01 ? ((x06 & ((~x03 & (x00 ? (x05 ? (x09 & (~x02 ^ x07) & (x04 ^ x10)) : ((~x02 & ~x04 & x07 & x09) | (x02 & x04 & ~x07 & ~x09 & ~x10))) : ((~x02 & ((~x07 & (x04 ? (~x10 & (x05 | (~x05 & x09))) : (x05 & x09))) | (~x04 & ~x05 & x07 & ~x09 & x10))) | (~x04 & x05 & ~x07 & ~x09 & x10)))) | (x07 & ((~x10 & (x02 ? (x03 & ((~x00 & (x04 ? x09 : (~x05 & ~x09))) | (~x05 & x09 & x00 & ~x04))) : (x05 & ((~x04 & ~x09) | (~x00 & x03 & x09))))) | (x00 & x02 & x03 & ((~x04 & x05 & ~x09 & x10) | (x04 & (x05 ? (x09 & x10) : ~x09)))))) | (x02 & x03 & ~x07 & ((~x00 & ~x09 & ((x05 & x10) | (x04 & ~x05 & ~x10))) | (x00 & x04 & ~x05 & x09 & x10))))) | (~x06 & (x09 ? (x00 ? (x04 ? (x02 ? (~x03 & (x05 ? (~x07 & x10) : (x07 & ~x10))) : (x03 & x07 & (~x05 ^ x10))) : ((x02 & x03 & ((x07 & ~x10) | (~x05 & ~x07 & x10))) | (~x02 & ~x03 & ~x05 & x07 & x10))) : (x10 & ((x03 & (x02 ? ((~x05 & x07) | (x04 & x05 & ~x07)) : (x04 & x07))) | (~x02 & ~x03 & x04 & ~x05 & ~x07)))) : ((~x07 & ((x00 & ((~x02 & ~x03 & ~x05 & x10) | (x02 & x03 & x04 & x05 & ~x10))) | (~x02 & ~x10 & ((~x03 & ~x04 & x05) | (~x00 & x03 & x04 & ~x05))))) | (x00 & ~x02 & ~x03 & x04 & x05 & x10)))) | (~x05 & x07 & ~x09 & ~x10 & x00 & x02 & x03 & ~x04)) : (x03 ? (x02 ? (x00 ? ((x10 & ((x05 & ((~x04 & x06 & x07 & x09) | (x04 & ~x09 & (x06 ^ ~x07)))) | (~x04 & ~x05 & (x06 ? ~x07 : (x07 & x09))))) | (~x09 & ~x10 & ((~x06 & x07 & ~x04 & x05) | (x06 & ~x07 & x04 & ~x05)))) : ((x09 & ((x04 & x06 & (x05 ? (x07 & ~x10) : (~x07 & x10))) | (~x06 & ~x10 & (~x05 ^ x07)))) | (~x05 & ~x06 & ~x09 & (x04 ? (x07 & ~x10) : (~x07 & x10))))) : ((~x09 & (x00 ? (x04 ? (x07 & (x05 ? (~x06 & x10) : (x06 & ~x10))) : (~x06 & ~x07 & (~x05 ^ x10))) : (x06 & ((~x05 & x07 & ~x10) | (~x04 & x10 & (~x07 | (~x05 & x07))))))) | (~x00 & x05 & ~x06 & x07 & x09 & x10))) : (x04 ? ((~x10 & (x00 ? ((x02 & x05 & ~x06 & x07) | (~x02 & ~x05 & ~x07 & x09)) : (~x09 & ((~x02 & (x07 ? ~x06 : ~x05)) | (x02 & x05 & x06 & ~x07))))) | (~x00 & x10 & (x02 ? ((~x05 & ~x06 & x09) | (x05 & x06 & x07 & ~x09)) : ((x05 & ~x06 & x07 & x09) | (~x05 & x06 & ~x07 & ~x09))))) : ((x02 & ((~x06 & x07 & ((x00 & (x05 ? (x09 & ~x10) : (~x09 & x10))) | (~x00 & ~x05 & x09 & ~x10))) | (~x05 & x06 & ((~x07 & ~x09 & ~x10) | (~x00 & x09 & x10))))) | (~x02 & ~x05 & x06 & x07 & x09 & x10)))))) | (x04 & ((x02 & (x03 ? (x07 ? ((~x00 & ~x01 & x06 & ((~x08 & ~x09 & ~x10) | (~x05 & x09 & x10))) | (x00 & x01 & ~x05 & ~x06 & ~x08 & ~x09 & x10)) : (x00 ? ((~x01 & ~x06 & ((x05 & x09 & ~x10) | (~x05 & ~x08 & ~x09 & x10))) | (x01 & x05 & ~x08 & ~x09 & ~x10)) : ((x01 & ((~x05 & ~x06 & ~x09 & x10) | (x05 & x06 & ~x08 & x09 & ~x10))) | (~x05 & x06 & ~x08 & ~x09 & ~x10)))) : (~x08 & (x05 ? (x07 & x10 & (x01 ? ((~x06 & ~x09) | (~x00 & (~x06 ^ ~x09))) : (x06 & ~x09))) : ((x09 & ((~x00 & x07 & (x01 ? (x06 & x10) : (~x06 & ~x10))) | (x00 & ~x01 & ~x06 & ~x07 & x10))) | (x00 & ~x07 & ~x09 & (x01 ? (~x06 & x10) : (x06 & ~x10)))))))) | (~x08 & ((~x03 & ((~x09 & ((~x00 & ((~x02 & ~x10 & ((x01 & (x05 ? ~x06 : (x06 & ~x07))) | (x06 & x07 & ~x01 & ~x05))) | (~x06 & ~x07 & x10 & ~x01 & ~x05))) | (x01 & ~x02 & x05 & x06 & x07 & (~x10 | (x00 & x10))))) | (x01 & ~x07 & x09 & ((~x06 & x10 & ~x00 & ~x05) | (x00 & ~x02 & (x05 ? (~x06 & x10) : (x06 & ~x10))))))) | (~x02 & x03 & ((x01 & (x00 ? (x10 & ((~x06 & ~x07 & ~x09) | (x05 & x06 & x07 & x09))) : (~x10 & ((~x05 & x06 & (x07 ^ x09)) | (x05 & ~x06 & ~x07 & x09))))) | (x00 & ~x01 & ~x07 & ((x05 & (x06 ? (x09 & ~x10) : (~x09 & x10))) | (~x05 & ~x06 & x09 & ~x10))))))) | (x00 & ~x01 & ~x02 & ~x03 & ~x05 & x06 & x07 & x09 & x10))) | (~x08 & ((~x04 & ((x01 & (x03 ? ((~x09 & ((~x06 & ((~x10 & ((~x02 & x05 & ~x07) | (x00 & (x02 ? (~x05 & ~x07) : (x05 & x07))))) | (~x00 & x10 & (x02 ? (x05 & x07) : ~x07)))) | (~x02 & ~x05 & x06 & x10 & (x00 | (~x00 & x07))))) | (~x07 & x09 & ((x00 & ((x02 & ~x05 & x06 & ~x10) | (~x02 & ~x06 & x10))) | (x02 & x05 & x06 & x10)))) : (x02 ? (x07 & ((~x00 & ~x06 & (x05 ? (x09 & ~x10) : (~x09 & x10))) | (x00 & ~x05 & x06 & ~x09 & ~x10))) : (x00 ? (~x07 & ~x09 & (x05 ? (x06 & x10) : (~x06 & ~x10))) : (x09 & ~x10 & (x05 ? ~x06 : (x06 & x07))))))) | (~x01 & (x00 ? ((x07 & (x03 ? (x05 & x10 & ((~x06 & x09) | (x02 & x06 & ~x09))) : ((x06 & (x02 ? (x05 ? (x09 & ~x10) : (~x09 & x10)) : (x09 & ~x10))) | (~x02 & ~x05 & ~x06 & x09 & x10)))) | (~x06 & x09 & ~x10 & ~x02 & ~x03 & x05)) : ((~x06 & ((~x07 & ((~x02 & x10 & ((x05 & ~x09) | (~x03 & ~x05 & x09))) | (x02 & ~x03 & x05 & x09 & ~x10))) | (x07 & x09 & ~x10 & ~x02 & ~x03 & ~x05))) | (x06 & ~x07 & x09 & ~x10 & ~x02 & ~x03 & ~x05)))) | (x00 & x02 & x03 & x05 & x06 & ~x07 & ~x09 & x10))) | (x01 & ~x02 & ~x05 & x07 & x10 & ((~x00 & x03 & ~x06 & x09) | (x00 & ~x03 & x06 & ~x09))))) | (~x00 & x01 & ~x02 & ~x03 & ~x04 & ~x05 & x06 & ~x07 & ~x09 & x10);
  assign z13 = (x03 & ((x02 & ((x01 & ((~x08 & (x00 ? ((~x06 & ((~x07 & ((x04 & ((~x09 & ~x10) | (~x05 & x09 & x10))) | (~x04 & x05 & ~x09 & ~x10))) | (~x04 & x07 & (x05 ? (x09 & x10) : ~x10)))) | (x04 & x05 & ((x06 & ~x09 & x10) | (~x07 & x09 & ~x10)))) : ((~x10 & ((x04 & ((x05 & x06 & x09) | (~x05 & ~x06 & x07 & ~x09))) | (~x04 & ~x05 & x06 & ~x07 & x09))) | (~x04 & x05 & x09 & x10 & (x06 ^ ~x07))))) | (x05 & ((x06 & ((x08 & ((x07 & ~x09 & (x00 ? (x04 ^ x10) : ~x04)) | (~x00 & ~x07 & x09 & (~x04 ^ x10)))) | (x00 & x04 & x07 & x09 & x10))) | (x00 & ~x04 & ~x06 & ~x07 & x08 & x09 & ~x10))) | (~x07 & x08 & ~x09 & x10 & ~x05 & x06 & x00 & x04))) | (~x01 & ((~x07 & (x00 ? (x04 ? (~x09 & ((x05 & (x06 ? (x08 & x10) : ~x10)) | (x08 & ~x10 & ~x05 & x06))) : ((x10 & ((~x06 & ~x08 & ~x09) | (~x05 & (x06 ? (~x08 & x09) : (x08 & ~x09))))) | (x05 & ~x06 & x08 & ~x09 & ~x10))) : (x08 ? ((x04 & ((~x05 & ~x06 & ~x09 & x10) | (x05 & ~x10 & (x06 | (~x06 & x09))))) | (~x05 & x06 & x09 & ~x10)) : ((~x04 & ~x05 & ~x06 & ~x09 & ~x10) | (x06 & x09 & x10 & x04 & x05))))) | (x08 & ((x07 & ((~x04 & ((x10 & ((~x00 & (x05 ? ~x06 : (x06 & x09))) | (x00 & x05 & x06 & x09))) | (~x00 & ~x05 & ~x06 & x09 & ~x10))) | (x00 & x04 & ((~x06 & x09 & ~x10) | (~x05 & (x06 ? (x09 & ~x10) : (~x09 & x10))))))) | (x06 & x09 & x10 & ~x00 & x04 & ~x05))))) | (~x05 & x10 & ((x00 & x07 & x09 & (x04 ? (x06 & ~x08) : (~x06 & x08))) | (~x07 & x08 & ~x09 & ~x00 & ~x04 & x06))))) | (~x02 & ((x01 & ((~x05 & ((x10 & (((x04 ? (x06 & ~x08) : (~x06 & x08)) & (x00 ? (~x07 & ~x09) : (x07 & x09))) | (~x07 & ~x08 & x09 & ~x00 & ~x04 & x06))) | (~x10 & ((x00 & ~x06 & x08 & (x04 ? ~x07 : (x07 & x09))) | (x07 & ~x08 & x09 & ~x00 & ~x04 & x06))) | (~x07 & ~x08 & x09 & ~x00 & x04 & x06))) | (x05 & (x09 ? ((~x04 & x07 & ((x00 & x08 & (~x06 ^ ~x10)) | (~x08 & ~x10 & ~x00 & ~x06))) | (~x00 & x04 & ~x06 & x08 & ~x10)) : ((~x00 & ((x06 & ((x04 & ((x08 & ~x10) | (~x07 & ~x08 & x10))) | (x08 & x10 & ~x04 & x07))) | (~x04 & ~x06 & x07 & (~x08 ^ ~x10)))) | (~x07 & ~x08 & ~x10 & x00 & ~x04 & x06)))) | (~x04 & ((~x06 & ~x07 & ~x08 & x09 & ~x10) | (x08 & ~x09 & x10 & x00 & x06 & x07))))) | (~x01 & (x08 ? (x04 ? ((x00 & x05 & x06 & ~x07 & x09) | (~x05 & ~x06 & x07 & ~x09 & x10)) : (~x10 & ((~x05 & (x00 ? (x09 & (x06 ^ ~x07)) : (~x09 & (~x07 | (~x06 & x07))))) | (x06 & ~x07 & x00 & x05)))) : ((~x06 & ((~x07 & (x00 ? ((~x04 & x05 & ~x09 & x10) | (x04 & ~x05 & x09 & ~x10)) : (~x09 & ((x04 & ~x05 & x10) | (x05 & ~x10))))) | (~x05 & x07 & x09 & x00 & ~x04))) | (~x00 & x06 & x07 & ((x04 & x09 & (~x05 ^ x10)) | (~x04 & ~x05 & ~x09 & x10)))))) | (~x07 & x08 & x10 & ((~x05 & x06 & x09 & x00 & ~x04) | (~x00 & x05 & ~x06 & ~x09))))) | (~x04 & ~x08 & x09 & ((~x00 & ~x01 & ((~x05 & ~x06 & x07 & x10) | (x05 & x06 & ~x07 & ~x10))) | (x06 & x07 & x10 & x00 & x01 & ~x05))))) | (x05 & ((~x07 & ((~x04 & (x06 ? ((x00 & ((~x01 & ~x03 & ((x02 & x08 & (~x09 ^ x10)) | (~x02 & ~x08 & x09 & x10))) | (x01 & ~x02 & x08 & ~x09 & x10))) | (~x01 & ~x02 & ~x03 & ~x08 & ~x09 & x10)) : ((x08 & ((~x03 & ((x00 & ~x01 & x09 & (~x10 | (~x02 & x10))) | (~x00 & x01 & x02 & ~x09 & x10))) | (~x00 & x01 & x02 & ~x09 & ~x10))) | (~x03 & ~x08 & ((~x01 & ~x02 & ((x09 & x10) | (x00 & ~x09 & ~x10))) | (x01 & x02 & ~x09 & ~x10)))))) | (~x03 & ((x00 & ((x04 & ((~x06 & ((x02 & x08 & (x01 ? ~x10 : (x09 & x10))) | (~x01 & ~x02 & ~x08 & (x09 ^ x10)))) | (~x01 & x06 & ~x10 & ((x08 & x09) | (~x02 & ~x08 & ~x09))))) | (x01 & ~x02 & x06 & x09 & (~x08 ^ x10)))) | (~x00 & ~x01 & ~x02 & x04 & x06 & x08 & ~x09))))) | (~x03 & ((x00 & ((x07 & ((~x02 & ((x04 & ((~x09 & ((x01 & (x10 ? x06 : x08)) | (x08 & ~x10 & ~x01 & x06))) | (~x01 & x06 & ~x08 & x09 & x10))) | (~x08 & ~x09 & ~x10 & ~x01 & ~x04 & x06))) | (~x01 & x02 & ~x04 & ~x10 & (x06 ? (~x08 & x09) : (x08 & ~x09))))) | (x01 & ~x02 & x04 & ~x06 & ~x08 & x09 & x10))) | (x07 & ((~x00 & ((x06 & ((x04 & ((x01 & x02 & x08 & ~x09 & x10) | (~x01 & ~x02 & ~x08 & x09 & ~x10))) | (~x09 & ((x01 & ~x10 & (x02 ^ x08)) | (~x01 & ~x02 & ~x04 & ~x08 & x10))) | (x08 & x09 & x10 & ~x01 & x02 & ~x04))) | (x04 & ((~x06 & x09 & ((x01 & (x02 ? (x08 & x10) : (~x08 & ~x10))) | (~x01 & x02 & x08 & ~x10))) | (~x01 & ~x02 & ~x08 & ~x09 & ~x10))))) | (x06 & x08 & ~x09 & x10 & ~x01 & x02 & ~x04))))))) | (~x05 & ((~x03 & ((~x04 & (x01 ? ((x06 & ((~x07 & ((x10 & ((x00 & (x02 ? x08 : (~x08 & x09))) | (~x00 & x02 & x08 & x09))) | (~x00 & ~x02 & ~x08 & x09 & ~x10))) | (x00 & x07 & x08 & ~x10 & (x02 ^ ~x09)))) | (x00 & ~x06 & ~x08 & ((x02 & x09 & (x07 ^ ~x10)) | (x07 & ~x09 & (~x10 | (~x02 & x10)))))) : (x00 ? (x02 & ((~x06 & ((~x08 & ~x09 & ~x10) | (~x07 & x08 & x09 & x10))) | (x06 & x07 & ~x08 & ~x09 & ~x10))) : ((x10 & ((~x02 & ((x06 & ~x08 & x09) | (~x06 & ~x07 & x08 & ~x09))) | (~x07 & ~x08 & x02 & x06))) | (x06 & x07 & ~x08 & x09 & ~x10))))) | (x04 & (x07 ? ((~x08 & ((x00 & ((~x01 & ~x02 & ~x06 & ~x09 & x10) | (x01 & x02 & x06 & x09 & ~x10))) | (~x00 & ~x01 & ~x02 & ~x06 & x09 & x10))) | (~x00 & ~x01 & x02 & x06 & x08 & ~x09 & ~x10)) : (x00 ? ((~x01 & ((x06 & ~x08 & x09 & x10) | (x02 & ~x06 & x08 & ~x09 & ~x10))) | (x08 & x09 & ~x10 & x01 & x02 & ~x06)) : ((~x10 & (x01 ? (~x02 & (x06 ? ~x08 : (x08 & ~x09))) : (x02 & (x06 ? (x08 & x09) : (~x08 & ~x09))))) | (x02 & x08 & x10 & (x01 ? (~x06 & x09) : (x06 & ~x09))))))) | (~x00 & ~x01 & ~x02 & x07 & x08 & (x06 ? (~x09 & x10) : (x09 & ~x10))))) | (~x00 & x01 & x06 & ~x07 & ~x09 & ((x02 & x04 & ~x08 & x10) | (~x02 & ~x04 & x08 & ~x10))))) | (~x06 & x07 & x08 & ~x09 & x10 & ~x00 & ~x01 & ~x03 & x04);
  assign z14 = (~x01 & ((x04 & ((((~x00 & ~x02 & x05 & ~x06 & x07) | (x00 & x02 & ~x05 & x06 & ~x07)) & ((x03 & x08 & ~x09 & x10) | (~x03 & ~x08 & x09 & ~x10))) | (x09 & (x02 ? (x00 ? ((x10 & (x03 ? ((~x05 & ~x06 & ~x07) | (x07 & x08 & x05 & x06)) : ((~x07 & ~x08 & x05 & ~x06) | (x07 & x08 & ~x05 & x06)))) | (~x06 & ~x07 & x08 & ~x03 & x05)) : (~x10 & (x03 ? ((~x05 & ~x06 & ~x08) | (~x07 & x08 & x05 & x06)) : (~x07 & ((~x06 & x08) | (x05 & x06 & ~x08)))))) : (~x08 & ((x06 & ((~x00 & x03 & ~x05 & x07 & x10) | (~x03 & (x00 ? (x05 & (x07 ^ ~x10)) : (~x05 & ~x10))))) | (~x06 & ~x07 & ~x10 & ~x00 & x03 & x05))))) | (~x09 & ((~x03 & (((x07 ? (x08 & ~x10) : (~x08 & x10)) & ((x00 & ~x02 & ~x05 & x06) | (x05 & ~x06 & ~x00 & x02))) | (~x02 & ((~x10 & ((x00 & ((x05 & x06 & ~x07) | (~x05 & ~x06 & x07 & ~x08))) | (~x00 & x05 & x06 & ~x07 & x08))) | (~x00 & ((~x05 & ~x06 & ~x07 & x10) | (x07 & ~x08 & x05 & x06))))) | (~x06 & x07 & x08 & x10 & (x00 ? x02 : ~x05)))) | (~x00 & ~x02 & x05 & ~x08 & ~x10 & ~x06 & ~x07))))) | (~x04 & ((x09 & (x10 ? (x00 ? (x03 & x05 & x08 & (x02 ? (~x07 | (~x06 & x07)) : (x06 & x07))) : (x02 ? ((~x06 & x07 & x08 & ~x03 & x05) | (x03 & x06 & (x05 ? (x07 & ~x08) : (~x07 & x08)))) : (~x07 & (x03 ? (~x05 & ~x06) : (x05 ? (~x06 & x08) : (x06 & ~x08)))))) : ((~x03 & ((x02 & (x00 ? ((~x07 & ~x08 & x05 & x06) | (x07 & x08 & ~x05 & ~x06)) : (x06 ? (x08 & (x05 ^ x07)) : (~x07 & ~x08)))) | (~x00 & x08 & ((x05 & ~x06 & x07) | (~x02 & x06 & ~x07))))) | (x07 & ((x03 & ((~x02 & (x00 ? (x05 ? (~x06 & x08) : ~x08) : (x06 & (x05 ^ x08)))) | (~x00 & x02 & ~x05 & ~x06 & ~x08))) | (x00 & ~x02 & x05 & x06 & ~x08)))))) | (~x09 & (x06 ? ((x08 & ((~x02 & ((x00 & x05 & (x03 ? (~x07 & ~x10) : (x07 & x10))) | (~x00 & x03 & ~x05 & ~x07 & ~x10))) | (~x00 & x02 & ~x03 & (x05 ? (x07 & ~x10) : (x07 ^ ~x10))))) | (~x00 & ~x02 & x03 & x10 & (x05 ? x07 : (~x07 & ~x08)))) : ((x03 & ((~x08 & ((x00 & ((~x02 & x05 & x07) | (x02 & ~x05 & ~x07 & ~x10))) | (x07 & x10 & ~x00 & ~x05))) | (~x02 & ~x05 & ~x07 & x08 & ~x10))) | (x00 & x02 & ~x03 & ((~x05 & (x07 ? (~x08 & ~x10) : (x08 & x10))) | (x05 & x07 & ~x08 & x10)))))) | (x08 & x10 & ~x06 & ~x07 & x00 & ~x02 & x03 & x05))) | (x03 & ((~x05 & ((x00 & x09 & x10 & ((~x06 & x07 & x08) | (~x07 & ~x08 & ~x02 & x06))) | (~x00 & ~x02 & x06 & x07 & ~x08 & ~x09 & ~x10))) | (x00 & x02 & x05 & ~x06 & ~x07 & ~x08 & ~x09 & x10))))) | (x01 & ((x09 & ((~x02 & ((x04 & (((x05 ^ ~x06) & ((x00 & ~x03 & ~x07 & ~x08 & x10) | (~x00 & x03 & x07 & x08 & ~x10))) | (~x00 & ((~x03 & x07 & ((~x06 & x08 & x10) | (~x08 & ~x10 & ~x05 & x06))) | (~x05 & x06 & ~x07 & x08 & ~x10))) | (x07 & x08 & ~x10 & x00 & ~x03 & ~x05))) | (x05 & ((~x06 & ((~x04 & ((x00 & ((~x07 & x08 & x10) | (~x03 & x07 & ~x10))) | (~x07 & x08 & x10 & ~x00 & x03))) | (~x00 & ~x07 & ~x08 & (~x03 ^ x10)))) | (x00 & x06 & ((~x03 & ((x07 & x08 & x10) | (~x08 & ~x10 & ~x04 & ~x07))) | (x07 & ~x08 & ~x10 & x03 & ~x04))))) | (~x04 & ~x05 & ((x00 & x06 & ((x03 & ~x10 & (~x07 ^ x08)) | (~x08 & x10 & ~x03 & ~x07))) | (~x00 & ~x03 & ~x06 & ~x07 & x08))))) | (x02 & (x04 ? (x00 ? ((x07 & ((~x06 & ((~x03 & x05 & ~x08) | (x10 & (x03 ? (~x05 ^ x08) : (~x05 & x08))))) | (x08 & ~x10 & x03 & x06))) | (x06 & x08 & x10 & (x03 ? x05 : (~x05 & ~x07)))) : ((x06 & ((~x03 & x07 & ~x08 & (x05 ^ x10)) | (x03 & ~x05 & ~x07 & x08 & ~x10))) | (~x07 & ~x08 & x10 & ~x03 & ~x06))) : (x00 ? ((x05 & ((~x03 & ~x10 & (x06 ? x07 : (~x07 & ~x08))) | (x03 & x06 & x07 & ~x08 & x10))) | (x03 & ~x05 & ~x06 & x08 & (x07 ^ ~x10))) : ((x07 & ~x08 & ((~x06 & ~x10 & ~x03 & x05) | (x03 & (x05 ? (~x06 & x10) : (x06 & ~x10))))) | (~x03 & ~x05 & x06 & x08 & x10))))) | (x08 & x10 & x06 & ~x07 & ~x04 & ~x05 & x00 & x03))) | (~x09 & (x10 ? ((~x02 & ((x04 & ((~x05 & (x00 ? ((~x03 & x07 & x08) | (~x07 & ~x08 & x03 & ~x06)) : (x06 & ~x08 & (x03 ^ ~x07)))) | (x06 & ~x07 & ~x08 & ~x00 & x03 & x05))) | (~x00 & ((~x03 & x05 & ((x06 & ~x07 & x08) | (~x04 & (x06 ? (x07 & ~x08) : ~x07)))) | (x03 & ~x04 & ~x05 & ~x06 & x08))))) | (x02 & ((x08 & ((x00 & ((x03 & x06 & x07 & (x04 | (~x04 & x05))) | (~x06 & ~x07 & ((~x04 & x05) | (~x03 & x04 & ~x05))))) | (~x00 & ~x03 & ~x04 & x05 & x06 & x07))) | (~x00 & ~x05 & ~x06 & x07 & ~x08 & (x03 ^ ~x04)))) | (~x00 & ~x03 & ~x04 & x07 & x08 & ~x05 & x06)) : (x02 ? ((x03 & ((~x08 & ((x00 & x07 & (x04 ? (~x05 & ~x06) : (x05 & x06))) | (~x00 & x04 & x05 & x06 & ~x07))) | (~x04 & ~x07 & x08 & (x05 ? x06 : ~x00)))) | (x06 & x07 & ~x08 & ~x00 & ~x04 & x05)) : (x00 ? (((x06 ? (~x07 & x08) : (x07 & ~x08)) & (x03 ? (~x04 & ~x05) : (x04 & x05))) | (x03 & ~x05 & x06 & ~x07 & ~x08)) : ((x05 & ((x03 & ((x07 & x08 & x04 & ~x06) | (~x07 & ~x08 & ~x04 & x06))) | (~x03 & ~x04 & ~x06 & x07 & ~x08))) | (~x03 & ~x05 & x06 & x07 & ~x08)))))) | (x00 & ~x02 & x03 & x04 & x05 & x06 & ~x07 & x08 & x10))) | (~x03 & ~x04 & x09 & ((x00 & ~x02 & ~x06 & ~x10 & (x05 ? (~x07 & ~x08) : (x07 & x08))) | (~x08 & x10 & x06 & ~x07 & ~x00 & x02 & x05)));
  assign z15 = (x04 & ((~x06 & (x10 ? ((x01 & ((x07 & (x00 ? ((x09 & ((x02 & (x03 ? (~x05 & ~x08) : (x05 & x08))) | (~x05 & x08 & ~x02 & ~x03))) | (~x02 & x03 & x05 & ~x08 & ~x09)) : ((~x05 & (x02 ? (x03 ? (x08 & ~x09) : (~x08 & x09)) : (x03 ? (x08 & x09) : (~x08 & ~x09)))) | (x02 & ~x03 & x05 & x08 & ~x09)))) | (~x05 & ~x07 & ((x02 & ((x00 & (x03 ? ~x09 : (~x08 & x09))) | (~x00 & ~x03 & x08 & x09))) | (~x00 & ~x02 & x03 & x08 & ~x09))))) | (~x01 & ((~x02 & (x00 ? ((x03 & x09 & (x08 ? x05 : x07)) | (~x03 & ~x05 & x07 & x08 & ~x09)) : ((~x03 & x07 & ~x08 & x09) | (x03 & x05 & ~x07 & x08 & ~x09)))) | (x00 & ((x03 & ((~x05 & ~x07 & ~x08 & ~x09) | (x02 & x07 & (x05 ? (x08 & x09) : (~x08 & ~x09))))) | (x02 & x05 & ((~x07 & ~x08 & x09) | (~x03 & x07 & x08 & ~x09))))))) | (x00 & ~x02 & x03 & ~x08 & ~x09 & x05 & ~x07)) : (x00 ? ((x02 & ((x09 & ((~x01 & ~x07 & x08 & (~x03 ^ ~x05)) | (x01 & x03 & x05 & x07 & ~x08))) | (~x03 & x05 & ~x09 & ((x07 & x08) | (~x01 & ~x07 & ~x08))))) | (~x01 & ~x02 & ((~x03 & ~x05 & (x07 ^ ~x09)) | (x03 & x05 & ~x07 & x09)))) : (x09 ? ((x01 & ((~x02 & ~x03 & (x05 ? (~x07 & x08) : (x07 & ~x08))) | (x02 & x03 & ~x05 & x07 & x08))) | (~x03 & x05 & ((~x01 & x07 & x08) | (~x02 & ~x07 & ~x08)))) : ((x07 & ((x05 & ((x01 & (x02 ? (~x03 & ~x08) : (x03 & x08))) | (~x01 & x02 & x03 & ~x08))) | (~x01 & ~x02 & ~x03 & ~x05 & x08))) | (x02 & x03 & ~x05 & ~x07 & (x01 ^ x08))))))) | (x06 & ((x01 & ((x03 & (x09 ? ((x08 & (x00 ? (x10 & (x02 ? (~x05 & x07) : (x05 & ~x07))) : (~x05 & ~x10 & (x02 ^ x07)))) | (x07 & ~x08 & x10 & ~x00 & x02 & x05)) : (x00 ? (~x08 & ~x10 & (x02 ? (~x05 & ~x07) : (x05 & x07))) : (x08 & ((~x02 & ~x05 & (~x07 | (x07 & x10))) | (x02 & x05 & ~x07 & x10)))))) | (~x03 & ((x07 & ((x08 & ((~x02 & ((~x00 & x09 & (x05 ^ x10)) | (x00 & ~x05 & ~x09 & x10))) | (x00 & x02 & (x05 ? (~x09 & x10) : (x09 & ~x10))))) | (x05 & ~x08 & x09 & (x00 ? ~x10 : (~x02 & x10))))) | (~x07 & x08 & ~x09 & x10 & x00 & ~x02 & x05))) | (~x07 & ~x08 & ~x09 & x10 & ~x00 & ~x02 & ~x05))) | (~x01 & ((x00 & (x05 ? (x09 & ((x02 & x10 & (x03 ? (~x07 & ~x08) : (x07 & x08))) | (~x02 & ~x03 & ~x07 & ~x08 & ~x10))) : ((x08 & ((x02 & ((~x09 & x10 & x03 & x07) | (~x03 & ~x07 & x09 & ~x10))) | (~x02 & ~x07 & ~x09 & ~x10))) | (~x08 & x09 & x10 & ~x02 & x03 & x07)))) | (~x00 & (x07 ? ((~x02 & ~x08 & ((x03 & x05 & x10) | (~x03 & ~x05 & ~x09 & ~x10))) | (x02 & ~x03 & x05 & x08 & ~x10)) : (x02 ? ((~x03 & ((x05 & x08 & x10) | (~x05 & ~x08 & x09 & ~x10))) | (x03 & x05 & ~x08 & x09)) : (~x09 & ((~x08 & x10 & x03 & ~x05) | (x08 & ~x10 & ~x03 & x05)))))) | (x02 & ~x03 & x05 & ~x07 & ~x08 & x09 & x10))) | (~x07 & x08 & ~x09 & x10 & x00 & x02 & ~x03 & ~x05))) | (x00 & ~x01 & ~x05 & x10 & ((x02 & ~x03 & x07 & ~x08 & x09) | (~x02 & x03 & ~x07 & x08 & ~x09))))) | (~x04 & ((~x00 & ((x03 & (x02 ? (x01 ? ((~x08 & ((~x10 & ((~x05 & ~x06 & x07 & ~x09) | (x05 & ((~x07 & ~x09) | (x06 & x07 & x09))))) | (~x05 & x06 & x07 & ~x09 & x10))) | (x08 & x09 & x10 & ~x05 & x06 & x07)) : ((~x07 & ((~x05 & ~x06 & x10 & (x08 ^ x09)) | (x05 & x08 & x09 & ~x10))) | (x06 & x07 & ((x08 & x09 & ~x10) | (x05 & (x08 ? (x09 & x10) : (~x09 & ~x10))))))) : ((x05 & ((x10 & ((x01 & ~x06 & ((~x07 & ~x08 & x09) | (x08 & ~x09))) | (~x01 & x06 & ~x07 & ~x08 & ~x09))) | (~x01 & x06 & x08 & ~x10 & (x07 ^ x09)))) | (~x01 & ((~x05 & ((~x06 & x07 & x08 & ~x09 & x10) | (x06 & ((~x07 & x08 & ~x09 & x10) | (x07 & ~x08 & x09 & ~x10))))) | (x06 & ~x07 & x08 & ~x09 & ~x10))) | (~x07 & x08 & x09 & ~x10 & x01 & ~x05 & x06)))) | (~x03 & (((~x02 ^ x06) & ((~x08 & x09 & x10 & ~x01 & x05 & x07) | (x08 & ~x09 & ~x10 & x01 & ~x05 & ~x07))) | (~x01 & ((~x07 & ((~x05 & ((x02 & (x06 ? (x09 & x10) : (~x08 & ~x10))) | (~x02 & ~x06 & ~x08 & x09 & x10))) | (~x08 & x09 & x10 & ~x02 & x05 & x06))) | (x02 & x05 & x08 & ((x06 & x09 & ~x10) | (~x06 & x07 & ~x09 & x10))))) | (x01 & ((x10 & ((x08 & ((x02 & (x05 ? (~x07 & x09) : (~x06 & x07))) | (x05 & x06 & x07 & ~x09) | (~x02 & ~x05 & ~x06 & ~x07 & x09))) | (~x07 & ~x08 & ~x09 & ~x02 & ~x05 & ~x06))) | (~x02 & ~x05 & x06 & ~x07 & ~x08 & x09))))) | (~x01 & ~x09 & ~x10 & ((~x06 & x07 & x08 & ~x02 & ~x05) | (x02 & x05 & x06 & ~x07 & ~x08))))) | (x00 & ((x08 & (x10 ? ((~x03 & ((x02 & ~x06 & (x01 ? (x07 & (x05 ^ x09)) : (x05 ? (~x07 & x09) : ~x09))) | (~x01 & ~x02 & x06 & ~x09 & (x05 ^ x07)))) | (x06 & ~x07 & ((~x01 & ~x02 & ((~x05 & ~x09) | (x03 & x05 & x09))) | (x02 & x03 & ~x05 & x09)))) : ((x03 & (x05 ? ((x06 & ((x01 & ((x07 & x09) | (~x02 & ~x07 & ~x09))) | (~x01 & x02 & x07 & x09))) | (x07 & x09 & ~x01 & ~x06)) : ((~x01 & ~x07 & ~x09 & (~x06 | (x02 & x06))) | (~x02 & ~x06 & x07 & x09)))) | (x01 & ~x02 & ((~x03 & x05 & ~x06 & ~x07 & x09) | (~x05 & x06 & x07 & ~x09))) | (x06 & ~x07 & ~x09 & ~x01 & ~x03 & ~x05)))) | (~x08 & (x03 ? ((~x02 & (x01 ? ((~x05 & x06 & x07 & x09 & x10) | (x05 & ~x06 & ~x07 & ~x09)) : (~x05 & x06 & ~x07 & (~x09 ^ x10)))) | (~x07 & ~x10 & ((~x01 & x05 & x06 & x09) | (x02 & ~x05 & ~x06 & ~x09)))) : ((x10 & ((~x02 & ((~x01 & ~x09 & (x05 ? (x06 & x07) : (~x06 & ~x07))) | (x01 & ~x05 & ~x06 & ~x07 & x09))) | (x01 & x02 & x07 & (x05 ? (x06 & x09) : ~x09)))) | (x05 & ~x06 & ~x10 & ((~x02 & ~x07 & x09) | (~x01 & x02 & x07 & ~x09)))))) | (x01 & ~x03 & ((x02 & x05 & ~x06 & ~x07 & ~x09 & x10) | (~x02 & ~x05 & x06 & x07 & x09 & ~x10))))) | (x01 & ~x02 & ~x03 & ~x05 & x06 & x07 & x08 & x09 & x10))) | (x02 & ~x07 & ((~x00 & ((x06 & x08 & ~x09 & x10 & x01 & ~x03 & x05) | (~x01 & x03 & ~x05 & ~x06 & ~x08 & x09 & ~x10))) | (x00 & x01 & ~x03 & x05 & ~x06 & ~x08 & ~x09 & ~x10)));
  assign z16 = (~x09 & ((~x00 & (x02 ? ((x03 & (x01 ? ((~x06 & ((~x04 & x07 & (x05 ? (x08 & x10) : ~x10)) | (~x07 & ~x08 & ~x10 & x04 & x05))) | (x04 & x06 & x08 & (x05 ? (x07 & x10) : (~x07 & ~x10)))) : ((x05 & ~x06 & ((~x07 & ~x08 & x10) | (x04 & x08 & (x07 ^ x10)))) | (~x04 & ~x05 & x06 & (x07 ? (x08 & x10) : (~x08 & ~x10)))))) | (~x03 & ((x07 & ((x10 & ((x01 & (x04 ? (x05 ? (~x06 & ~x08) : (x06 & x08)) : (x05 ? (x06 & ~x08) : ~x06))) | (~x01 & x04 & ~x05 & x06 & ~x08))) | (~x01 & x06 & ~x10 & (~x05 ^ x08)))) | (x01 & ~x07 & ~x10 & ((x06 & x08 & x04 & x05) | (~x04 & ~x05 & ~x08))))) | (~x08 & x10 & ~x06 & ~x07 & x01 & ~x04 & ~x05)) : ((x01 & (x03 ? ((x08 & ((x04 & ((x05 & x06 & ~x07) | (~x05 & ~x06 & x07 & x10))) | (~x04 & ~x05 & ~x06 & x07 & ~x10))) | (~x04 & ((x06 & ~x07 & (x05 ? ~x10 : (~x08 & x10))) | (~x08 & x10 & ~x06 & x07)))) : ((x05 & ((~x04 & ((~x08 & x10 & x06 & ~x07) | (x08 & ~x10 & ~x06 & x07))) | (x04 & ~x06 & x07 & x08 & x10))) | (x04 & ~x05 & ((x08 & ~x10 & ~x06 & ~x07) | (x06 & x07 & (~x08 ^ ~x10))))))) | (x10 & ((x05 & ((~x01 & ~x04 & ~x06 & x08 & (x03 ^ x07)) | (x03 & x04 & x06 & x07 & ~x08))) | (~x01 & ~x03 & ~x05 & ((~x07 & (x04 ? (~x06 ^ x08) : (x06 & ~x08))) | (x07 & x08 & ~x04 & x06))))) | (~x05 & ~x06 & x07 & ~x08 & ~x01 & ~x03 & ~x04)))) | (x00 & ((x04 & (x07 ? (x01 ? ((~x03 & ((x05 & x06 & ~x08 & x10) | (~x02 & ~x05 & ~x06 & x08 & ~x10))) | (~x08 & ((~x02 & ((x05 & ~x06 & x10) | (x03 & x06 & (x05 ^ x10)))) | (x02 & x03 & x05 & ~x06 & ~x10)))) : (x05 ? ((~x02 & ((x03 & x08 & x10) | (~x08 & ~x10 & ~x03 & x06))) | (~x08 & ~x10 & ~x03 & ~x06)) : ((x02 & ~x06 & x10 & (~x03 ^ x08)) | (x06 & x08 & ~x02 & x03)))) : ((x01 & ((~x06 & ((~x02 & ~x03 & x08 & (x05 | (~x05 & x10))) | (~x08 & ~x10 & x02 & x03))) | (x02 & x03 & ((x05 & (~x08 ^ ~x10)) | (~x08 & x10 & ~x05 & x06))))) | (~x05 & ~x06 & x08 & ((x02 & x03 & x10) | (~x01 & ~x02 & ~x03 & ~x10)))))) | (~x08 & ((~x04 & ((~x02 & ((x05 & ~x07 & (x01 ? (x10 & (~x03 ^ x06)) : (~x06 & ~x10))) | (~x01 & ~x05 & x07 & ~x10 & (x03 ^ x06)))) | (x01 & x02 & x05 & ((x03 & x07 & (~x06 ^ ~x10)) | (~x07 & x10 & ~x03 & x06))))) | (~x05 & ~x06 & ~x07 & x10 & ~x01 & ~x02 & x03))) | (~x03 & x08 & ((~x04 & (x01 ? ((x02 & ((x05 & x06 & ~x07 & ~x10) | (~x05 & x10 & (x06 ^ ~x07)))) | (~x02 & ~x05 & ~x06 & x07 & x10)) : ((x06 & ~x07 & x10 & ~x02 & x05) | (x02 & ~x05 & ~x06 & x07 & ~x10)))) | (x06 & ~x07 & x10 & ~x01 & x02 & ~x05))))) | (~x01 & ~x02 & ~x03 & x05 & ~x06 & x10 & (x04 ? (x07 & ~x08) : (~x07 & x08))))) | (x09 & ((x02 & ((x01 & (x03 ? (x10 ? ((x00 & x08 & ((x05 & ~x06 & x07) | (x04 & ~x05 & ~x07))) | (~x06 & x07 & ~x08 & ~x00 & x04 & ~x05)) : ((~x04 & x07 & ((x00 & ~x08 & (x05 ^ x06)) | (~x06 & x08 & ~x00 & x05))) | (~x00 & x04 & ~x07 & (x05 ? (x06 & x08) : (~x06 & ~x08))))) : ((~x10 & ((~x00 & ~x05 & (x04 ? (x06 ? (~x07 & ~x08) : (x07 & x08)) : (~x06 & ~x08))) | (x06 & ~x07 & ~x08 & x00 & ~x04 & x05))) | (x00 & x05 & x06 & ~x08 & x10 & (x04 ^ x07))))) | (x05 & ((~x01 & ((~x07 & ((~x04 & ((~x06 & ((~x00 & x08 & (x03 ^ x10)) | (~x08 & ~x10 & x00 & ~x03))) | (x00 & x06 & x10 & (~x08 | (x03 & x08))))) | (x00 & ~x03 & x04 & x08 & ~x10))) | (x04 & ~x06 & x07 & ~x08 & ((~x03 & x10) | (x00 & x03 & ~x10))))) | (x08 & x10 & x06 & x07 & x00 & x03 & x04))) | (~x01 & ~x05 & ((~x07 & (x00 ? ((~x03 & x04 & ~x06 & x08 & x10) | (~x08 & ~x10 & x03 & ~x04)) : (x08 & (x03 ? (x10 ? ~x04 : x06) : (x04 ? (x06 & x10) : ~x10))))) | (~x00 & x04 & x06 & x07 & (x08 ? x03 : ~x10)))))) | (~x02 & (x07 ? (x06 ? ((x04 & (x00 ? ((~x01 & ((x08 & x10 & ~x03 & x05) | (~x08 & ~x10 & x03 & ~x05))) | (~x05 & x08 & x01 & x03)) : (x01 & ((x03 & (x05 ? (x08 & x10) : (~x08 & ~x10))) | (~x08 & ~x10 & ~x03 & x05))))) | (~x00 & ~x04 & ((~x01 & ~x03 & ~x05 & (~x08 ^ ~x10)) | (x05 & ~x08 & ~x10 & x01 & x03)))) : ((x05 & ((x08 & (x00 ? ((x01 & x03 & ~x04) | (x04 & ~x10 & ~x01 & ~x03)) : (x10 & (x01 ? (x03 & ~x04) : (~x03 & x04))))) | (x00 & x01 & ~x03 & x04 & ~x08 & x10))) | (~x04 & ~x05 & ~x08 & x10 & x00 & x01 & x03))) : (x04 ? (x06 ? ((~x00 & x03 & ~x08 & ((~x05 & ~x10) | (~x01 & x05 & x10))) | (x00 & ~x01 & ~x03 & ~x05 & x08 & ~x10)) : ((x05 & ((x00 & ((~x03 & ~x08 & ~x10) | (x08 & x10 & x01 & x03))) | (~x00 & ~x01 & x03 & x08 & x10))) | (~x00 & x01 & ~x03 & ~x05 & ~x08 & x10))) : ((~x08 & ((x00 & x10 & (x01 ? (~x05 & ~x06) : (x03 & x05))) | (~x00 & x01 & x03 & x05 & ~x06))) | (~x00 & x01 & ~x03 & x08 & ~x10 & x05 & ~x06))))) | (~x05 & ~x10 & ((x00 & ((~x06 & x07 & x08 & ~x01 & ~x03 & x04) | (x06 & ~x07 & ~x08 & x01 & x03 & ~x04))) | (~x00 & x01 & x03 & x07 & ~x08 & ~x04 & x06))))) | (x03 & ~x05 & ((x00 & ~x07 & ~x10 & ((~x01 & x02 & x04 & x06 & x08) | (x01 & ~x02 & ~x04 & ~x06 & ~x08))) | (~x08 & x10 & ~x06 & x07 & ~x02 & x04 & ~x00 & ~x01)));
  assign z17 = (x05 & ((x06 & ((x00 & (x03 ? ((x07 & (x01 ? (x02 & ((~x09 & x10 & x04 & x08) | (~x04 & ~x08 & x09 & ~x10))) : ((~x04 & ((x08 & ~x09 & ~x10) | (~x02 & (x08 ? x09 : (~x09 & x10))))) | (x04 & ~x08 & x09 & ~x10)))) | (~x10 & ((x04 & ~x07 & (x01 ? (x02 ? (x08 & ~x09) : x09) : (x02 ? (x08 & x09) : (~x08 & ~x09)))) | (x01 & ~x02 & ~x04 & x08 & ~x09)))) : (x04 ? (x07 & (x01 ? (~x08 & (x02 ? (x09 & ~x10) : (~x09 & x10))) : (x08 & ~x09 & (x02 | (~x02 & x10))))) : (x01 ? (x07 & x10 & (x02 ? (x08 & x09) : (x08 ^ x09))) : ((~x09 & ((~x07 & ~x08 & x10) | (~x02 & (x08 ? ~x07 : ~x10)))) | (~x02 & x07 & x08 & x09 & x10)))))) | (x04 & ((~x00 & (x03 ? ((~x07 & x10 & ((~x01 & x09 & (x02 ^ ~x08)) | (x01 & ~x02 & x08 & ~x09))) | (~x02 & x07 & ~x08 & ~x09 & ~x10)) : ((~x10 & ((~x09 & ((x01 & (x08 ? x07 : x02)) | (~x01 & ~x02 & ~x07 & x08))) | (~x01 & x02 & x07 & ~x08 & x09))) | (x01 & x02 & ~x07 & x10 & (x08 ^ ~x09))))) | (~x01 & x02 & x03 & x07 & ~x08 & x09 & x10))) | (~x04 & ((~x00 & ~x02 & ((~x07 & ((~x08 & ((x01 & ~x09 & (x03 ^ x10)) | (~x01 & x03 & x09 & ~x10))) | (~x01 & x03 & x08 & ~x09))) | (~x01 & x07 & x08 & (x03 ? (x09 & x10) : (~x09 & ~x10))))) | (x01 & x02 & ~x03 & ~x07 & x08 & ~x09 & x10))))) | (~x06 & ((~x07 & ((~x01 & ((((x02 & ~x08 & ~x09 & x10) | (~x02 & x08 & x09 & ~x10)) & (x00 ? (x03 & ~x04) : (~x03 & x04))) | (~x09 & ((~x00 & x03 & ((x02 & x04 & x08) | (~x02 & ~x04 & ~x08 & x10))) | (x00 & ~x02 & ~x03 & x08 & x10))) | (x00 & ~x04 & x09 & (x02 ? (x08 & ~x10) : (~x08 & x10))))) | (x04 & ((x01 & x02 & ((x00 & ~x03 & x09 & (~x08 ^ ~x10)) | (~x09 & ((x03 & x08 & x10) | (~x00 & ~x08 & ~x10))))) | (x08 & x09 & x10 & ~x00 & ~x02 & x03))) | (x01 & ~x03 & (x00 ? ((~x02 & ~x04 & x08 & x09 & x10) | (x02 & ~x08 & ~x09 & ~x10)) : (~x04 & ((x02 & ~x08 & x09 & x10) | (~x02 & x08 & ~x09 & ~x10))))))) | (x07 & (x04 ? ((~x01 & ((x00 & ~x10 & ((x02 & ~x03 & ~x08 & x09) | (~x02 & x03 & x08 & ~x09))) | (~x08 & x09 & x10 & ~x00 & ~x02 & ~x03))) | (~x00 & x01 & x02 & x09 & x10 & ~x03 & x08)) : (x01 ? ((x00 & x03 & ((~x02 & ~x08 & x09 & x10) | (x02 & x08 & ~x09 & ~x10))) | (x08 & ((~x00 & ~x10 & (x02 ? ~x09 : (~x03 & x09))) | (~x02 & ~x03 & ~x09 & x10)))) : (x09 & ((~x00 & x02 & ~x03 & (~x08 ^ x10)) | (x00 & ~x02 & ~x08 & ~x10)))))) | (x00 & ~x01 & ~x02 & x03 & x04 & ~x08 & x09 & x10))) | (~x04 & ((~x00 & ~x01 & ~x10 & ((x02 & x03 & ~x07 & x08 & x09) | (~x02 & ~x03 & x07 & ~x08 & ~x09))) | (x07 & ~x08 & x09 & x10 & x00 & x01 & x02 & ~x03))))) | (~x05 & ((~x07 & (x10 ? ((x00 & ((~x02 & ((~x01 & ((~x03 & x04 & ~x06 & ~x08 & x09) | (x03 & ~x04 & x06 & x08 & ~x09))) | (x06 & x08 & x09 & x01 & ~x03 & ~x04))) | (x01 & ((x02 & ((x03 & ((x04 & ~x08 & x09) | (~x04 & ~x06 & x08 & ~x09))) | (~x03 & x04 & x06 & ~x08 & x09))) | (x03 & ~x04 & ~x06 & ~x08 & x09))))) | (x08 & ((~x00 & ~x03 & ~x06 & ((x01 & ~x04 & (~x09 | (~x02 & x09))) | (~x01 & ~x02 & x04 & ~x09))) | (x04 & x06 & x09 & ~x01 & ~x02 & x03))) | (~x00 & x01 & x02 & ~x08 & ((~x03 & x04 & ~x06 & x09) | (x03 & ~x04 & x06 & ~x09)))) : ((~x00 & (x03 ? ((~x09 & ((~x01 & (x02 ? (~x06 & x08) : (x04 & x06))) | (x01 & ~x02 & ~x06 & x08))) | (x01 & x02 & x04 & x09 & (~x08 | (x06 & x08)))) : ((~x08 & ((~x01 & ~x04 & (x02 ? (x06 & x09) : (~x06 & ~x09))) | (x01 & x02 & x04 & x06 & x09))) | (x01 & x04 & ~x06 & x08 & (~x09 | (x02 & x09)))))) | (x00 & (x01 ? ((~x02 & ((x03 & x04 & ~x06 & x08 & x09) | (~x03 & ~x04 & x06 & ~x08 & ~x09))) | (x03 & ~x04 & ~x09 & (~x06 ^ x08))) : ((x02 & ((~x03 & x06 & x08 & x09) | (~x04 & ~x06 & ~x08 & ~x09))) | (~x02 & ~x03 & x04 & x06 & x09)))) | (~x01 & ~x02 & x03 & x04 & ~x06 & ~x08 & x09)))) | (x07 & ((~x06 & (x10 ? (x03 ? ((x01 & ((x08 & ((x00 & x09 & (x02 ^ x04)) | (~x00 & x02 & ~x04 & ~x09))) | (~x00 & x04 & ~x08 & (x02 ^ ~x09)))) | (~x00 & ~x01 & ~x02 & ~x04 & ~x08 & ~x09)) : ((~x09 & ((x02 & ((x00 & x08 & (~x01 ^ x04)) | (~x00 & x01 & x04 & ~x08))) | (~x02 & ~x04 & ~x08 & x00 & ~x01))) | (~x00 & x04 & x09 & ((~x02 & (~x08 | (x01 & x08))) | (~x01 & x02 & x08))))) : (x01 ? ((x08 & ((x00 & ((~x02 & x03 & ~x04 & ~x09) | (x02 & x09))) | (~x00 & ~x02 & ~x03 & ~x04 & ~x09))) | (~x00 & ~x02 & ~x03 & x04 & ~x08 & ~x09)) : (x04 & ~x08 & ((x00 & x02 & x03 & x09) | (~x02 & ~x03 & ~x09)))))) | (x06 & (x01 ? (~x02 & ~x09 & ((~x00 & (x03 ? (~x04 & ~x10) : (x10 & (x04 | (~x04 & x08))))) | (~x04 & ~x08 & x10 & x00 & ~x03))) : (x04 ? ((~x09 & ((~x00 & x02 & ~x03 & (~x08 ^ x10)) | (~x02 & ((x00 & ((~x08 & ~x10) | (x03 & x08 & x10))) | (~x08 & x10 & ~x00 & x03))))) | (x00 & ~x02 & ~x03 & x08 & x09)) : (x09 & ((~x00 & ~x03 & (x02 ? (x08 & x10) : (~x08 & ~x10))) | (x00 & ~x02 & x03 & ~x08 & x10)))))) | (x00 & x01 & x02 & ~x03 & ~x04 & ~x08 & ~x09 & x10))) | (x06 & x09 & ((~x00 & ~x01 & ~x02 & ~x08 & x10 & x03 & ~x04) | (x00 & x01 & x02 & x08 & ~x10 & ~x03 & x04))))) | (x00 & ((~x08 & ((~x07 & (x01 ? (x02 & ~x03 & ((~x04 & x06 & ~x09 & x10) | (x04 & ~x06 & x09 & ~x10))) : (~x02 & x03 & ~x04 & ~x09 & (~x06 ^ ~x10)))) | (~x02 & x03 & x07 & x09 & x10 & (x01 ? (x04 & x06) : (~x04 & ~x06))))) | (x04 & x06 & ~x07 & x08 & ~x10 & ((~x01 & ~x02 & x03 & x09) | (x01 & x02 & ~x03 & ~x09))))) | (~x00 & x01 & x02 & x03 & ~x04 & ~x06 & x07 & x08 & x09 & ~x10);
  assign z18 = (x03 & ((x07 & (x10 ? ((~x04 & (x06 ? (x08 ? ((~x01 & ((~x09 & (x00 ? (~x02 ^ ~x05) : ~x05)) | (~x00 & ~x02 & x05 & x09))) | (x00 & x01 & (x02 ? (x05 & ~x09) : (~x05 & x09)))) : ((~x00 & ~x09 & ((x02 & ~x05) | (x01 & ~x02 & x05))) | (~x01 & ~x02 & ~x05 & x09))) : ((x02 & ((x00 & ~x08 & (x01 ? (~x05 & x09) : (x05 & ~x09))) | (~x05 & x08 & (x09 ? ~x01 : ~x00)))) | (x01 & ~x02 & x05 & ~x08 & (~x09 | (x00 & x09)))))) | (x01 & x04 & ((~x09 & ((~x05 & (x00 ? (x02 ? x08 : (~x06 & ~x08)) : (~x02 & x06))) | (~x00 & ~x02 & x05 & x06 & x08))) | (~x00 & x05 & x09 & (x02 ? (~x06 ^ x08) : (~x06 & x08)))))) : ((x06 & (x01 ? ((x04 & x08 & ((x00 & ((~x05 & ~x09) | (x02 & x05 & x09))) | (~x00 & ~x02 & ~x05 & x09))) | (~x00 & ~x02 & ~x04 & ~x05 & x09)) : (x02 ? ((~x04 & ((~x00 & x09 & (~x05 ^ x08)) | (x00 & x05 & ~x08 & ~x09))) | (x00 & x04 & (x05 ? x08 : (~x08 & ~x09)))) : ((~x09 & (x00 ? (x04 ^ ~x05) : (x04 & ~x05))) | (~x05 & x08 & x09 & x00 & ~x04))))) | (~x06 & ((x09 & ((~x01 & ((x05 & ~x08 & (x00 ? (x02 ^ x04) : (x02 & x04))) | (~x00 & ~x02 & ~x04 & ~x05 & x08))) | (~x00 & x01 & x02 & x04 & x05 & x08))) | (x01 & x02 & ~x09 & ((~x00 & (x04 ? ~x05 : (x05 & x08))) | (~x05 & ~x08 & x00 & ~x04))))) | (~x00 & x01 & x02 & ~x04 & x05 & ~x08 & x09)))) | (~x07 & ((~x10 & (x02 ? (x00 ? ((x05 & ((~x04 & ((x01 & ~x06 & (~x09 | (x08 & x09))) | (~x01 & x06 & x08 & x09))) | (~x08 & ~x09 & ~x01 & x04))) | (~x01 & ~x05 & x09 & ((x06 & x08) | (x04 & ~x06 & ~x08)))) : (x01 ? (~x05 & (x04 ? (x06 & x08) : (~x06 & ~x09))) : (x05 & x06 & ~x08 & (~x04 ^ ~x09)))) : (x09 ? ((x01 & ((x00 & ((~x04 & x06 & ~x08) | (~x06 & x08 & x04 & ~x05))) | (x05 & ((x04 & x06 & x08) | (~x06 & ~x08 & ~x00 & ~x04))))) | (~x00 & ~x01 & ~x04 & (x05 ? (~x06 & x08) : ~x08))) : ((~x05 & ((~x00 & ((~x04 & x06 & ~x08) | (x01 & x04 & ~x06 & x08))) | (x06 & x08 & x00 & ~x04))) | (x05 & x06 & ~x08 & ~x00 & ~x01 & ~x04))))) | (x10 & ((x08 & ((x02 & ((x04 & ~x09 & ((~x00 & ~x06 & (x01 ^ x05)) | (x05 & x06 & x00 & x01))) | (~x05 & x06 & x09 & ~x00 & ~x01 & ~x04))) | (x00 & ((~x02 & x05 & ((~x04 & x06 & x09) | (x01 & ((x04 & x06 & x09) | (~x06 & ~x09))))) | (~x01 & ~x04 & ~x05 & x06 & ~x09))))) | (~x02 & ~x08 & ((~x01 & ((~x04 & ((x00 & (x05 ? (x06 & ~x09) : (~x06 & x09))) | (~x00 & ~x05 & x06 & ~x09))) | (~x00 & x04 & ~x05 & ~x06 & x09))) | (~x05 & x06 & x09 & x00 & x01 & ~x04))))) | (~x01 & ~x05 & ((~x06 & x08 & x09 & ~x00 & ~x02 & x04) | (x00 & x02 & ~x04 & x06 & ~x08 & ~x09))))) | (~x02 & x04 & ~x00 & x01 & x05 & ~x06 & x08 & ~x09 & x10))) | (~x03 & (x06 ? ((x02 & (x05 ? (x00 ? ((~x04 & ((~x07 & x10 & (x01 ? (x08 ^ ~x09) : (x08 & ~x09))) | (x08 & ~x10 & ~x01 & x07))) | (x01 & x04 & ((~x07 & ~x08 & x09 & ~x10) | (x07 & x08 & ~x09 & x10)))) : (x10 & ((~x01 & x04 & x09 & (~x07 ^ x08)) | (~x07 & x08 & ~x09 & x01 & ~x04)))) : ((x07 & ((~x08 & ((x00 & ~x10 & (x01 ? (x04 & x09) : (~x04 & ~x09))) | (~x04 & x09 & x10 & (~x01 | (~x00 & x01))))) | (~x00 & x01 & ~x04 & x08 & x09 & ~x10))) | (~x00 & x01 & ~x04 & ~x07 & x08 & ~x09 & ~x10)))) | (~x02 & (x00 ? ((~x08 & ((x01 & ~x04 & ((~x05 & x07 & x09 & x10) | (~x09 & ~x10 & x05 & ~x07))) | (x07 & ~x09 & ~x10 & ~x01 & x04 & ~x05))) | (x04 & x08 & ((~x01 & ((~x09 & ~x10 & x05 & ~x07) | (~x05 & (x07 ? (~x09 & x10) : (x09 & ~x10))))) | (~x05 & ~x07 & ~x09 & ~x10)))) : (x01 ? (x04 ? (~x07 & ~x08 & (x05 ? (~x09 & ~x10) : (x09 & x10))) : (x07 & x08 & x10 & (x05 ^ x09))) : ((~x05 & x07 & x08 & ~x09 & ~x10) | (~x07 & ((x04 & ~x08 & (x05 ? (~x09 & x10) : (x09 & ~x10))) | (~x04 & x05 & x08 & x09 & ~x10))))))) | (~x07 & ~x08 & x09 & ~x10 & x00 & x01 & x04 & ~x05)) : (x01 ? (x04 ? ((~x00 & ((x10 & ((x02 & ((x05 & x07 & x08 & x09) | (~x05 & ~x07 & ~x09))) | (~x02 & x05 & ~x07 & ~x08 & x09))) | (~x02 & ((x05 & ~x09 & (x07 ? ~x08 : (x08 & ~x10))) | (~x05 & ~x07 & x08 & x09 & ~x10))))) | (x10 & ((~x02 & ((x05 & x07 & x08 & x09) | (x00 & ((x05 & ~x07 & x08) | (x07 & ~x08 & x09))))) | (~x07 & x08 & x09 & x00 & x02 & x05)))) : ((x02 & ((x08 & ((~x00 & (x05 ? (~x07 & ~x09) : (x07 & ~x10))) | (x00 & x05 & ~x07 & ~x09 & x10))) | (x00 & ~x08 & ~x10 & (x05 ? (x07 & ~x09) : (~x07 & x09))))) | (~x07 & ~x08 & x09 & ~x10 & x00 & ~x02 & x05))) : (x10 ? (x02 ? ((x07 & ((x05 & ((x09 & (x00 ? (~x08 | (x04 & x08)) : (~x04 & x08))) | (~x00 & x04 & x08 & ~x09))) | (x00 & ~x04 & ~x05 & ~x08 & ~x09))) | (~x07 & x08 & x09 & ~x00 & ~x04 & ~x05)) : (((x08 ^ ~x09) & ((~x05 & x07 & ~x00 & ~x04) | (x05 & ~x07 & x00 & x04))) | (~x04 & ~x05 & ~x07 & x08 & x09) | (x07 & ~x08 & ~x09 & ~x00 & x04 & x05))) : (x08 ? ((x05 & ((~x00 & ((~x04 & ~x07 & ~x09) | (~x02 & x04 & x09))) | (x00 & x02 & x04 & x09))) | (x02 & x04 & ~x05 & x07 & ~x09)) : (x00 ? ((~x09 & (x02 ? (x04 ? (x05 & x07) : (~x05 & ~x07)) : (~x04 & x05))) | (~x02 & ~x04 & x05 & x07 & x09)) : ((x02 & ~x05 & (x04 ? ~x09 : (~x07 & x09))) | (~x02 & x04 & ~x07 & x09)))))))) | (~x00 & x02 & ~x08 & ((~x01 & ~x05 & ((x04 & x06 & ~x07 & x09 & x10) | (~x04 & ~x06 & x07 & ~x09 & ~x10))) | (x01 & ~x04 & x05 & x06 & ~x07 & x09 & ~x10)));
  assign z19 = (~x03 & ((x01 & ((x07 & (x09 ? ((x04 & ((~x10 & ((~x00 & x02 & ~x05 & ~x06 & ~x08) | (~x02 & ((x05 & ~x06 & x08) | (x00 & (x05 ? x06 : (~x06 & ~x08))))))) | (~x00 & x02 & x06 & x10 & (~x05 ^ x08)))) | (x05 & ((~x00 & ~x04 & ~x06 & (x02 ? ~x10 : (~x08 & x10))) | (x00 & x02 & x06 & ~x08 & x10))) | (~x00 & ~x02 & ~x04 & ~x05 & ~x06 & ~x08 & ~x10)) : (x10 ? ((x02 & ((x08 & (x00 ? (x04 ? (x05 & ~x06) : (~x05 & x06)) : (x04 & ~x06))) | (~x00 & x05 & ~x08 & (~x04 | (x04 & x06))))) | (~x00 & ~x02 & ~x04 & x05 & ~x06 & x08)) : (x00 ? ((~x02 & x06 & (x08 ? x04 : ~x05)) | (~x04 & ~x05 & ~x06 & x08)) : ((x02 & ((~x04 & ~x05 & x06 & x08) | (~x06 & ~x08 & x04 & x05))) | (~x02 & ~x04 & x05 & ~x06 & ~x08)))))) | (~x07 & (x02 ? (x04 ? ((x09 & ((~x08 & x10 & ~x05 & x06) | (x05 & ((x00 & (x06 ? (~x08 & ~x10) : (x08 & x10))) | (~x08 & x10 & ~x00 & ~x06))))) | (x08 & ~x09 & ~x10 & ~x00 & ~x05 & x06)) : (x06 & x08 & ((x00 & ~x10 & (x05 ^ ~x09)) | (~x00 & ~x05 & ~x09 & x10)))) : ((~x08 & (x00 ? (x04 & ((x05 & ~x06 & x09 & ~x10) | (~x05 & x06 & ~x09 & x10))) : ((~x05 & ~x06 & x10 & (~x09 | (~x04 & x09))) | (x05 & x06 & x09 & ~x10)))) | (~x00 & x08 & ((~x04 & x05 & ~x06 & x09 & ~x10) | (~x09 & ((x04 & (x05 ? (~x06 & ~x10) : (x06 & x10))) | (~x04 & ~x05 & x06 & ~x10)))))))) | (x00 & ~x02 & x04 & ~x05 & x06 & x08 & x09 & ~x10))) | (~x01 & (x08 ? ((~x04 & ((~x09 & ((~x02 & (x07 ? (x00 ? (x10 & (x05 ^ ~x06)) : (x05 & x06)) : (x05 ? (~x06 & x10) : (x06 & ~x10)))) | (~x00 & x02 & ~x07 & (x05 ? (~x06 & x10) : (x06 & ~x10))))) | (x00 & x09 & ((x02 & ~x05 & x06 & (x07 ^ x10)) | (~x06 & x07 & x10 & ~x02 & x05))))) | (x02 & ~x09 & (x00 ? (x04 & ((~x05 & (x06 ? (~x07 & ~x10) : (x07 & x10))) | (x05 & x06 & ~x07 & x10))) : ((x07 & ~x10 & x05 & ~x06) | (x06 & x10 & x04 & ~x05))))) : (x07 ? (x02 ? ((x06 & ((x00 & ((x09 & x10 & x04 & x05) | (~x04 & ~x05 & ~x09 & ~x10))) | (~x00 & x04 & x05 & x09 & ~x10))) | (~x04 & ~x05 & ~x06 & ~x09 & (~x10 | (~x00 & x10)))) : ((x00 & ((x05 & x06 & ~x09 & ~x10) | (x04 & ~x05 & x09 & (~x06 ^ ~x10)))) | (~x06 & x09 & x10 & ~x00 & ~x04 & ~x05))) : (x00 ? (x06 & ((~x09 & ((x02 & (x04 ? ~x10 : (~x05 & x10))) | (~x02 & ~x04 & x05 & x10))) | (~x02 & ~x04 & ~x05 & x09 & x10))) : ((~x02 & ((x04 & x05 & ~x06 & ~x09 & x10) | (~x04 & ~x05 & x09 & ~x10))) | (x09 & ((x06 & ~x10 & x04 & x05) | (x02 & ~x06 & (x04 ? (~x05 & x10) : (x05 & ~x10))))) | (x02 & x05 & x06 & ~x09 & x10)))))) | (~x00 & ((~x07 & ((x02 & ~x09 & ((~x04 & ~x05 & ~x06 & x08 & x10) | (x06 & ~x08 & ~x10 & x04 & x05))) | (~x02 & x04 & ~x05 & x06 & x08 & x09 & ~x10))) | (x07 & ~x08 & x09 & ~x10 & x05 & x06 & ~x02 & ~x04))) | (x00 & ~x02 & ~x04 & x05 & x06 & ~x07 & x08 & x09 & ~x10))) | (x03 & ((x01 & (x10 ? (x00 ? ((x07 & (x05 ? (x02 ? (x08 & (x04 ? (~x06 & x09) : (x06 & ~x09))) : (~x08 & ((x06 & ~x09) | (~x04 & ~x06 & x09)))) : ((x02 & ~x08 & (x04 ? ~x06 : (x06 & ~x09))) | (~x02 & x04 & ~x06 & x08 & x09)))) | (x05 & ~x07 & ((x02 & x08 & (x04 ? (x06 & ~x09) : (~x06 & x09))) | (~x02 & x04 & ~x06 & ~x08 & ~x09)))) : ((x02 & ((x06 & ((x08 & ((~x05 & (x04 ? (x07 ^ ~x09) : (x07 & ~x09))) | (~x04 & x05 & ~x07 & x09))) | (~x04 & x05 & x07 & ~x08 & x09))) | (~x05 & ~x06 & x09 & ((x07 & ~x08) | (x04 & ~x07 & x08))))) | (~x06 & ~x07 & x08 & x09 & ~x02 & ~x04 & ~x05))) : (x04 ? ((~x02 & ((x07 & ((~x09 & (x05 ? (x00 ? (~x06 ^ x08) : (x06 | (~x06 & x08))) : (x06 & ~x08))) | (x00 & ~x05 & x06 & ~x08 & x09))) | (~x07 & ~x08 & x09 & ~x00 & ~x05 & x06))) | (~x00 & x02 & ((x05 & ~x07 & ~x09 & (~x08 | (~x06 & x08))) | (~x05 & ~x06 & x07 & x08 & x09)))) : (x02 ? ((~x05 & ((~x00 & ((x06 & ~x08 & x09) | (~x06 & x07 & x08 & ~x09))) | (x00 & ~x06 & ~x07 & ~x08 & x09))) | (x00 & x05 & x06 & ~x08 & (x07 ^ x09))) : (x08 & ((~x06 & (x00 ? (~x05 & x07) : ((~x07 & ~x09) | (x05 & x07 & x09)))) | (x00 & x06 & ~x07 & (x05 ^ ~x09)))))))) | (~x01 & (x08 ? ((x02 & (x05 ? ((x00 & ~x06 & ((~x04 & (x07 ? (~x09 & x10) : (x09 & ~x10))) | (x04 & x07 & ~x09 & ~x10))) | (~x07 & ~x09 & x10 & ~x00 & ~x04 & x06)) : ((x04 & ((x06 & ((x00 & ~x09 & (x07 ^ x10)) | (x09 & ~x10 & ~x00 & x07))) | (~x06 & ~x07 & x09 & x10))) | (x07 & x09 & ~x10 & ~x00 & ~x06)))) | (~x02 & (x04 ? ((x06 & ((x10 & ((x00 & ~x09 & (x05 ^ x07)) | (~x00 & ~x05 & x07 & x09))) | (~x00 & x05 & x09 & ~x10))) | (~x07 & x09 & ~x10 & ~x00 & ~x05 & ~x06)) : ((x05 & ~x06 & x07 & x09 & ~x10) | (~x09 & ((~x00 & ((~x06 & x07 & x10) | (x05 & x06 & ~x07 & ~x10))) | (~x06 & ~x07 & x10 & x00 & x05)))))) | (x00 & ~x04 & x05 & x06 & ~x07 & x09 & x10)) : (x06 ? ((~x07 & (x00 ? ((x02 & x04 & ~x05 & x09 & x10) | (~x02 & ~x04 & x05 & ~x09 & ~x10)) : (~x05 & x10 & (x02 ? (~x04 & x09) : (x04 & ~x09))))) | (~x00 & ~x02 & ~x04 & x05 & x09 & x10)) : ((x05 & ((~x04 & ((~x00 & ~x09 & (x02 ? (x07 & ~x10) : (~x07 & x10))) | (x09 & x10 & x00 & ~x07))) | (x00 & x02 & x04 & (x07 ? (x09 & x10) : ~x09)))) | (~x04 & ~x05 & ((~x00 & ~x10 & (x02 ? x09 : (x07 & ~x09))) | (x00 & ~x02 & x07 & x09 & x10))))))) | (~x00 & ~x02 & x04 & x06 & ~x09 & ((x05 & x07 & ~x08 & x10) | (~x05 & ~x07 & x08 & ~x10))))) | (x09 & ((x00 & ((x01 & x07 & ~x10 & ((x02 & x04 & x05 & ~x06 & x08) | (~x02 & ~x04 & ~x05 & x06 & ~x08))) | (~x08 & x10 & x06 & ~x07 & ~x01 & x02 & ~x04 & x05))) | (~x00 & x01 & x02 & ~x04 & ~x05 & ~x06 & x07 & x08 & x10)));
  assign z20 = (x09 & ((x01 & ((x00 & ((x06 & (x02 ? (x03 ? (x07 & ((x08 & (x04 ? (~x05 ^ x10) : (~x05 & x10))) | (~x08 & x10 & ~x04 & x05))) : ((x05 & ((~x07 & ~x08 & x10) | (~x04 & x07 & x08))) | (~x07 & ~x10 & x04 & ~x05))) : ((~x05 & ((~x03 & ~x08 & (x04 ? (x07 & x10) : (~x07 & ~x10))) | (~x07 & x08 & x03 & x04))) | (x03 & x05 & ((x08 & x10 & ~x04 & x07) | (~x08 & ~x10 & x04 & ~x07)))))) | (~x06 & (x02 ? (x03 & ~x08 & (x04 ? (~x10 & (x05 ^ x07)) : (x07 & x10))) : ((x04 & ((~x03 & ((x05 & x07 & ~x08 & x10) | (~x05 & ~x07 & x08 & ~x10))) | (x03 & ~x05 & x07 & ~x08 & x10))) | (x03 & ~x05 & ((x07 & ~x08 & ~x10) | (~x04 & ~x07 & x10)))))) | (x02 & ~x03 & x04 & x08 & ~x10 & x05 & ~x07))) | (~x00 & (x02 ? ((~x05 & ((x10 & ((x03 & ((x07 & x08 & x04 & ~x06) | (~x07 & ~x08 & ~x04 & x06))) | (~x03 & x04 & x06 & x07 & ~x08))) | (~x03 & ~x04 & ~x06 & x07 & x08 & ~x10))) | (x04 & x05 & ((x03 & x06 & ~x07 & (~x08 ^ x10)) | (x07 & x08 & x10 & ~x03 & ~x06)))) : ((x10 & ((x05 & ((~x03 & ~x04 & ~x06 & x07 & ~x08) | (x03 & x06 & (x04 ? (x07 & ~x08) : (~x07 & x08))))) | (~x03 & x08 & ((x04 & x06 & ~x07) | (~x05 & ~x06 & x07))) | (x03 & x04 & ~x05 & x06 & ~x07 & ~x08))) | (x05 & ~x10 & ((~x03 & ((x07 & x08 & ~x04 & ~x06) | (~x07 & ~x08 & x04 & x06))) | (x03 & x04 & x06 & ~x07 & x08)))))) | (~x03 & ~x04 & x07 & ((~x02 & ~x05 & ~x06 & x08 & ~x10) | (x02 & x05 & x06 & ~x08 & x10))))) | (~x01 & (x00 ? (x05 ? (x02 ? ((x03 & ((~x07 & ((x04 & (x06 ? (~x08 & x10) : (x08 & ~x10))) | (x08 & x10 & ~x04 & x06))) | (~x04 & x07 & (x06 ? (x08 & ~x10) : (~x08 & x10))))) | (x07 & ~x08 & ~x10 & ~x03 & ~x04 & ~x06)) : ((~x06 & ((x07 & ((~x03 & x10 & (x04 ^ ~x08)) | (~x08 & ~x10 & x03 & x04))) | (~x07 & x08 & x10 & ~x03 & ~x04))) | (~x03 & ~x04 & x06 & ~x08 & (x07 ^ x10)))) : ((x07 & ((~x06 & ((x02 & ~x08 & (x03 ? ~x10 : (~x04 & x10))) | (~x02 & ~x03 & ~x04 & x08 & x10))) | (~x02 & x06 & ((x04 & x08 & (x03 ^ x10)) | (x03 & ~x04 & (~x10 | (~x08 & x10))))))) | (~x03 & ~x04 & ~x07 & ~x08 & (x02 ? ~x10 : (~x06 & x10))))) : (x02 ? ((x06 & ((~x03 & ~x07 & ((~x04 & x05 & ~x08) | (x08 & ~x10 & x04 & ~x05))) | (x07 & ~x08 & x10 & x03 & x04 & x05))) | (~x04 & ~x06 & ((~x07 & (x03 ? (~x08 & (~x05 ^ x10)) : (x08 & x10))) | (~x03 & ~x05 & x07 & x08 & x10)))) : ((~x10 & ((~x07 & ((x03 & ((x04 & ~x06 & ~x08) | (x05 & x06 & x08))) | (~x06 & x08 & ~x03 & ~x04))) | (~x03 & x06 & x07 & (x04 ? (~x05 & ~x08) : (x05 & x08))))) | (~x06 & x10 & ((x07 & ~x08 & ~x04 & ~x05) | (~x03 & x04 & (x05 ? x07 : ~x08)))))))) | (~x02 & ~x03 & ((x00 & x05 & ((~x04 & x06 & x07 & x08 & x10) | (x04 & ~x06 & ~x07 & ~x08 & ~x10))) | (x08 & x10 & x06 & x07 & ~x00 & ~x04 & ~x05))) | (x00 & x02 & x03 & ~x04 & x05 & ~x06 & x07 & x08 & ~x10))) | (~x10 & ((~x09 & ((~x00 & (x05 ? ((~x06 & ((x02 & ((x03 & ((x01 & (x04 ? (x07 & x08) : (~x07 & ~x08))) | (x07 & ~x08 & ~x01 & ~x04))) | (~x01 & ~x03 & x04 & x07 & ~x08))) | (~x01 & ~x02 & ~x03 & x04 & ~x07 & ~x08))) | (~x04 & x07 & ~x08 & x01 & x02 & ~x03)) : (x03 ? ((x02 & (((~x08 | (~x04 & x08)) & (x01 ? (x06 & ~x07) : (~x06 & x07))) | (x06 & x07 & ~x01 & ~x04))) | (~x01 & ((~x02 & ((~x07 & x08 & ~x04 & ~x06) | (x07 & ~x08 & x04 & x06))) | (~x07 & x08 & x04 & x06)))) : ((x04 & ((~x06 & ((~x01 & ~x02 & ~x07 & x08) | (x01 & x07 & (~x08 | (~x02 & x08))))) | (~x01 & x02 & x06 & x07 & ~x08))) | (x01 & ~x02 & ~x04 & x06 & ~x08))))) | (~x02 & ((x00 & ((~x05 & (x01 ? ((x03 & x04 & ~x06 & ~x07 & x08) | (~x03 & ~x04 & x06 & x07 & ~x08)) : (~x03 & ~x07 & (x04 ? (x06 & ~x08) : (~x06 ^ x08))))) | (~x01 & x05 & ((x03 & x06 & (x04 ? (x07 & ~x08) : (~x07 & x08))) | (~x03 & ~x04 & ~x06 & ~x07 & x08))))) | (x03 & ~x05 & ~x06 & x07 & ~x08 & (~x01 ^ x04)))) | (x00 & ((~x01 & ((x06 & x07 & x08 & ((x03 & ~x04 & ~x05) | (x02 & (x03 ? (x04 & ~x05) : (~x04 & x05))))) | (~x07 & ~x08 & x05 & ~x06 & x02 & ~x03 & x04))) | (x01 & x02 & ~x03 & ~x07 & x08 & x04 & x06))))) | (~x02 & x08 & ((~x00 & x01 & ((~x03 & ~x04 & ~x05 & x06 & x07) | (x03 & x04 & x05 & ~x06 & ~x07))) | (x00 & ~x01 & x03 & ~x06 & x07 & x04 & x05))))) | (~x09 & ((x10 & (x00 ? (x01 ? ((x06 & ((x08 & (x04 ? (x07 & ((~x03 & ~x05) | (~x02 & x03 & x05))) : (~x07 & (x02 ? (x03 ^ ~x05) : (x03 & ~x05))))) | (x02 & x05 & ~x08 & (x03 ? x07 : ~x04)))) | (~x04 & x05 & ~x06 & ~x07 & (x02 ? ~x08 : (~x03 & x08)))) : ((x07 & ((x02 & ~x08 & ((~x03 & ~x04 & ~x05) | (x05 & x06 & x03 & x04))) | (~x03 & x04 & x05 & ~x06 & x08))) | (x06 & ~x07 & x08 & ~x02 & ~x03 & x04))) : (x04 ? (x06 ? ((x02 & ((x03 & x07 & (x01 ? (x05 ^ x08) : (~x05 & ~x08))) | (~x01 & ~x03 & x05 & ~x07 & ~x08))) | (~x03 & x05 & (x01 ? (~x07 & x08) : (~x02 & x07)))) : ((~x08 & (x01 ? (~x07 & (x02 ? (~x03 & x05) : (x03 & ~x05))) : (~x02 & x07 & (~x03 | (x03 & x05))))) | (~x05 & x07 & x08 & ~x01 & x02 & ~x03))) : ((~x07 & ((~x08 & (((x02 ? (~x03 & ~x05) : (x03 & x05)) & (x01 ^ ~x06)) | (x01 & ~x02 & ~x03 & x05 & ~x06))) | (~x01 & x08 & ((x02 & x06 & (x03 ^ ~x05)) | (~x05 & ~x06 & ~x02 & ~x03))))) | (x07 & x08 & x05 & x06 & ~x01 & x02 & ~x03))))) | (~x01 & x07 & x08 & ((~x04 & x05 & x06 & ~x00 & ~x02 & x03) | (x04 & ~x05 & ~x06 & x00 & x02 & ~x03))))) | (~x00 & x01 & x02 & x03 & ~x04 & x05 & ~x06 & x07 & ~x08 & x10);
  assign z21 = (~x02 & ((~x06 & ((~x05 & (x08 ? ((x04 & ((~x09 & ((x00 & ~x01 & (x03 ? (x07 & x10) : ~x07)) | (x01 & ~x07 & ((x03 & ~x10) | (~x00 & ~x03 & x10))))) | (x07 & x09 & x10 & ~x00 & x01 & x03))) | (x00 & ~x03 & ~x04 & ((x09 & ~x10 & x01 & x07) | (~x01 & (x07 ? (~x09 & ~x10) : (x09 & x10)))))) : (x10 ? ((x01 & ((~x09 & ((x00 & (x03 ? (~x04 & x07) : x04)) | (~x00 & ~x03 & ~x04 & ~x07))) | (~x00 & ~x03 & x04 & ~x07 & x09))) | (~x00 & ~x01 & x03 & x07 & ~x09)) : ((~x04 & ((x00 & (x01 ? (x03 & ~x09) : (x07 & x09))) | (~x00 & x01 & x07 & x09))) | (~x00 & x04 & ~x07 & x09 & (~x03 | (~x01 & x03))) | (x00 & ~x01 & x03 & x07 & ~x09))))) | (~x00 & (x03 ? (x05 & ~x07 & ((x08 & ((x01 & ~x09 & (x04 ^ x10)) | (x09 & x10 & ~x01 & ~x04))) | (~x01 & ~x04 & ~x08 & ~x09 & x10))) : ((x05 & x08 & (x01 ? ((x04 & x07 & ~x09 & ~x10) | (x09 & x10 & ~x04 & ~x07)) : (~x07 & x09 & (~x04 ^ x10)))) | (~x08 & ~x09 & x10 & ~x01 & x04 & x07)))) | (x00 & ((x05 & ((~x08 & ((x09 & ((x04 & ((x01 & x03 & (x07 ^ x10)) | (~x07 & ~x10 & ~x01 & ~x03))) | (~x04 & ~x07 & x10 & ~x01 & ~x03))) | (~x01 & ~x04 & x07 & ~x09 & ~x10))) | (x04 & x08 & x09 & ((x03 & x07 & x10) | (x01 & ~x03 & ~x10))))) | (~x07 & x08 & x09 & x01 & x03 & ~x04))) | (x07 & x08 & x09 & x10 & ~x04 & x05 & x01 & x03))) | (x06 & (x07 ? (x10 ? (x03 ? (x00 ? (~x04 & (x01 ? (x05 ? (x08 & ~x09) : (~x08 & x09)) : (x08 & (~x05 | (x05 & x09))))) : ((x01 & ~x08 & x09 & (x04 ^ x05)) | (~x01 & x04 & x05 & x08 & ~x09))) : ((~x00 & ((x05 & ((~x08 & ~x09 & ~x01 & x04) | (x01 & (x04 ? (x08 & x09) : (~x08 & ~x09))))) | (~x01 & x04 & ~x05 & x08 & ~x09))) | (~x05 & ~x08 & ~x09 & x00 & x01 & x04))) : ((~x03 & ((x05 & ((~x00 & ((~x01 & x08 & ~x09) | (~x08 & x09 & x01 & ~x04))) | (x00 & x01 & ~x04 & ~x09))) | (x00 & x04 & ~x05 & (x01 ? (x08 ^ x09) : ~x08)))) | (x00 & x01 & ((x08 & x09 & x04 & x05) | (x03 & ~x05 & ~x08 & ~x09))))) : ((x08 & (x01 ? ((x00 & ~x04 & x05 & (x03 ? (x09 & x10) : (~x09 & ~x10))) | (~x00 & x03 & x04 & ~x09 & x10)) : ((~x05 & ((x09 & (x00 ? ((~x04 & ~x10) | (~x03 & x04 & x10)) : ((~x04 & x10) | (~x03 & x04 & ~x10)))) | (x04 & ~x09 & ~x10 & x00 & x03))) | (~x04 & x05 & x10 & x00 & x03)))) | (x01 & x03 & ~x08 & ((~x10 & ((~x00 & x09 & (x04 ^ ~x05)) | (x05 & ~x09 & x00 & x04))) | (~x00 & ~x04 & ~x05 & ~x09 & x10)))))) | (x00 & x01 & ~x07 & x08 & ~x09 & x10 & (x03 ? (~x04 & ~x05) : (x04 & x05))))) | (x02 & ((x05 & ((x03 & (x04 ? (x00 ? ((x01 & ((~x06 & x09 & (x07 ? (x08 & ~x10) : (~x10 | (x08 & x10)))) | (x06 & ~x07 & ~x08 & ~x09 & x10))) | (~x08 & x09 & x10 & ~x01 & ~x06 & ~x07)) : ((~x10 & ((x01 & ((~x07 & ~x08 & ~x09) | (x06 & x07 & x08 & x09))) | (~x06 & ~x07 & ~x08 & x09))) | (~x01 & x07 & x08 & (x06 ? ~x09 : (x09 & x10))))) : ((~x09 & ((~x08 & ((x00 & ((x01 & x06 & ~x07) | (x07 & x10 & ~x01 & ~x06))) | (~x00 & x01 & ~x06 & x07 & x10))) | (~x01 & ((~x10 & ((x00 & (x06 ? (~x07 & x08) : x07)) | (x07 & x08 & ~x00 & ~x06))) | (~x07 & x08 & x10 & ~x00 & ~x06))))) | (~x07 & x08 & x09 & ~x10 & x00 & x01 & x06)))) | (~x03 & (x10 ? ((~x04 & (x01 ? (x06 & ((~x00 & ((~x07 & ~x08 & x09) | (x08 & ~x09))) | (x08 & x09 & x00 & ~x07))) : (x00 ? ((~x06 & ~x07 & x08 & ~x09) | (x06 & x07 & ~x08 & x09)) : (~x06 & (x07 ? (~x08 & x09) : ~x09))))) | (~x00 & x04 & ((~x01 & ~x07 & (x06 ? (x08 & ~x09) : (~x08 & x09))) | (x08 & ~x09 & x01 & ~x06)))) : ((~x08 & ((~x04 & (x00 ? ((~x07 & x09 & x01 & ~x06) | (~x01 & x06 & x07 & ~x09)) : (x01 & ((~x07 & ~x09) | (~x06 & x07 & x09))))) | (~x06 & x07 & ~x09 & x00 & x04))) | (x07 & x08 & x09 & x00 & ~x01 & ~x06)))) | (x00 & x01 & ~x06 & x07 & ~x08 & ~x09 & x10))) | (~x05 & (x08 ? ((x09 & ((x07 & ((~x03 & ((x04 & ((x00 & x10 & (x01 | (~x01 & x06))) | (~x00 & x01 & ~x06 & ~x10))) | (~x00 & ~x01 & ~x04 & ~x06 & ~x10))) | (x00 & x03 & ~x04 & (x01 ? (~x06 & x10) : (x06 & ~x10))))) | (~x01 & ~x06 & ~x07 & ((x04 & x10 & ~x00 & ~x03) | (~x04 & ~x10 & x00 & x03))))) | (~x03 & x06 & x07 & ((x00 & ~x10 & (x01 ? (~x04 & ~x09) : x04)) | (~x00 & x01 & ~x04 & ~x09 & x10)))) : (x10 ? ((~x01 & (x00 ? (x03 & (x04 ? (~x07 & ~x09) : (x06 & x09))) : (~x03 & ~x06 & x09 & (~x04 ^ x07)))) | (x06 & x07 & x09 & x00 & ~x03 & ~x04)) : (x00 ? ((x07 & ((x01 & ((x03 & x04 & ~x06 & x09) | (~x04 & x06 & ~x09))) | (x03 & ~x04 & x06 & x09))) | (x01 & ~x03 & x04 & ~x07 & x09)) : ((~x09 & ((~x03 & ((~x01 & (x04 ? (~x06 & ~x07) : (x06 & x07))) | (x01 & x04 & x06 & x07))) | (x01 & ((x04 & ~x06 & x07) | (x03 & ~x04 & x06 & ~x07))))) | (x06 & ~x07 & x09 & ~x01 & ~x03 & ~x04)))))) | (x00 & ~x01 & ~x03 & x04 & ~x06 & x07 & ~x08 & x09 & ~x10))) | (~x03 & ((x01 & ~x05 & ((x04 & ~x06 & ((~x00 & ~x07 & ~x10 & (x08 ^ ~x09)) | (x08 & ~x09 & x10 & x00 & x07))) | (x00 & ~x04 & x06 & ((x07 & x08 & x09 & x10) | (~x07 & ~x08 & ~x09 & ~x10))))) | (~x00 & ~x01 & ~x04 & x05 & x06 & x07 & x08 & ~x09 & x10)));
  assign z22 = (x07 & ((x02 & ((x06 & ((x01 & ((x08 & (x03 ? ((~x10 & ((x00 & ~x05 & (~x04 ^ x09)) | (~x00 & x04 & x05 & x09))) | (~x00 & x05 & ~x09 & (~x04 | (x04 & x10)))) : (x05 & ((~x04 & ~x09 & x10) | (~x00 & (~x04 ^ ~x09)))))) | (x05 & ~x10 & ((x00 & ~x08 & x09 & (~x03 ^ ~x04)) | (~x00 & x03 & x04 & ~x09))))) | (~x09 & ((~x04 & ((x10 & ((x00 & ((x03 & x05 & ~x08) | (~x05 & x08 & ~x01 & ~x03))) | (~x00 & ~x01 & ~x03 & x05 & ~x08))) | (~x08 & ~x10 & x03 & x05))) | (~x00 & ~x01 & x05 & ((~x03 & x08 & ~x10) | (~x08 & x10 & x03 & x04))))) | (~x00 & ~x01 & ~x03 & x04 & ~x05 & ~x08 & x09 & ~x10))) | (~x06 & (x00 ? ((~x04 & (x01 ? ((x03 & ((x05 & x08 & ~x10) | (~x05 & ~x08 & x09 & x10))) | (~x03 & ~x05 & ~x08 & x09 & ~x10)) : ((x10 & (x03 ? (~x09 & (~x05 ^ x08)) : (x09 & (x05 ^ x08)))) | (x03 & x05 & ~x08 & x09 & ~x10)))) | (~x01 & ((~x10 & ((x03 & ((x04 & x05 & x08) | (~x05 & ~x08 & x09))) | (~x03 & x04 & ~x05 & x08 & x09))) | (~x03 & x04 & x10 & (x05 ? (x08 & ~x09) : (~x08 & x09)))))) : (~x04 & ((~x01 & ((~x03 & ~x05 & ~x08 & x09 & ~x10) | (x05 & ((~x03 & ~x08 & ~x09 & ~x10) | (x03 & (x08 ? (x09 & ~x10) : (~x09 & x10))))))) | (~x08 & x09 & x10 & x01 & ~x03 & ~x05))))) | (x00 & ~x01 & x03 & x04 & x05 & ~x08 & x09 & x10))) | (~x02 & ((x00 & ((x04 & ((~x01 & ((~x03 & ((~x05 & x06 & ~x08 & ~x09 & x10) | (x05 & ~x06 & x08 & x09 & ~x10))) | (~x05 & ~x09 & ((x06 & x08 & ~x10) | (~x08 & x10 & x03 & ~x06))))) | (x03 & x06 & ((x05 & ((~x08 & x09 & ~x10) | (x01 & (x08 ? (x09 ^ x10) : (x09 & x10))))) | (x01 & ~x05 & x08 & x09 & x10))))) | (~x04 & ((x08 & (x06 ? ((~x01 & x03 & x05 & ~x09) | (x01 & x10 & ((~x05 & ~x09) | (~x03 & x05 & x09)))) : ((~x03 & ~x05 & ~x09 & ~x10) | (~x01 & ((~x03 & x09 & ~x10) | (x03 & ~x05 & ~x09 & x10)))))) | (~x03 & ~x05 & ~x06 & ~x08 & x09 & x10))) | (x01 & x03 & ~x05 & ~x06 & ~x08 & x09 & ~x10))) | (~x01 & ((x06 & ((~x00 & ((x08 & ((x10 & ((x03 & (x04 ? (~x05 & x09) : (x05 & ~x09))) | (~x03 & ~x04 & ~x05 & ~x09))) | (~x03 & x04 & x05 & ~x09 & ~x10))) | (x03 & ~x04 & ~x05 & ~x08 & ~x09 & x10))) | (x08 & x09 & ~x10 & ~x03 & ~x04 & x05))) | (~x00 & x03 & ~x06 & ~x08 & ~x09 & (x04 ? (~x05 ^ x10) : (x05 & ~x10))))) | (~x00 & ((x05 & ((x03 & ((x01 & ~x04 & ~x08 & x09 & x10) | (x04 & ~x06 & x08 & ~x09 & ~x10))) | (x01 & ~x03 & ~x06 & (x04 ? (x08 & x09) : ((~x09 & x10) | (~x08 & x09 & ~x10)))))) | (x01 & ~x04 & ~x05 & x10 & ((x03 & ~x06 & x08 & x09) | (~x03 & x06 & ~x08 & ~x09))))) | (x01 & x03 & ~x05 & ~x06 & ~x09 & (x04 ? (x08 & x10) : (~x08 & ~x10))))) | (x01 & ((~x05 & (x00 ? (~x03 & ((~x04 & ~x06 & x08 & x09 & x10) | (x04 & x06 & ~x08 & ~x09 & ~x10))) : (x03 & ~x06 & ((x04 & ~x08 & x09 & x10) | (~x04 & x08 & ~x09 & ~x10))))) | (~x06 & x08 & ~x09 & ~x10 & x00 & ~x03 & x04 & x05))))) | (~x07 & ((x01 & (x00 ? (x05 ? ((x09 & ((x10 & ((x03 & ((x02 & (x04 ? (~x06 & x08) : (x06 & ~x08))) | (~x04 & x08 & (~x06 | (~x02 & x06))))) | (x04 & ~x06 & x08 & ~x02 & ~x03))) | (x06 & ~x08 & ~x10 & ~x02 & ~x03 & x04))) | (x02 & ~x04 & x08 & ~x09 & ((x06 & ~x10) | (~x03 & ~x06 & x10)))) : (x02 ? (x10 ? ((~x03 & x04 & x06 & ~x08 & x09) | (x03 & ~x04 & x08 & (~x09 | (x06 & x09)))) : ((~x03 & x08 & (x04 ? (x06 & x09) : (~x06 & ~x09))) | (x03 & x04 & ~x06 & ~x08 & x09))) : ((~x08 & ((x03 & ((x04 & ~x06 & ~x09 & x10) | (~x04 & x06 & x09 & ~x10))) | (~x04 & x09 & ((~x06 & ~x10) | (~x03 & x06 & x10))))) | (x08 & ~x09 & ~x10 & ~x03 & x04 & x06)))) : (x04 ? (x05 ? ((x09 & ((x02 & ((~x08 & x10 & x03 & x06) | (x08 & ~x10 & ~x03 & ~x06))) | (~x02 & ~x03 & ~x06 & ~x10))) | (~x02 & ~x06 & ~x09 & x10 & (x03 ^ x08))) : ((~x02 & ~x08 & ~x10 & ((~x06 & x09) | (x03 & x06 & ~x09))) | (x02 & ~x03 & x06 & ~x09 & x10))) : ((~x03 & ((x05 & ((x02 & ~x08 & ~x09 & (~x06 ^ ~x10)) | (x08 & x09 & (x06 ? ~x02 : ~x10)))) | (~x05 & x06 & ~x08 & x09 & ~x10))) | (~x02 & x03 & x05 & ~x06 & ~x08 & x09 & ~x10))))) | (~x01 & (x00 ? (x03 ? ((x10 & ((x02 & ~x06 & ((x04 & ~x05 & (x08 ^ x09)) | (~x04 & x05 & ~x08 & ~x09))) | (~x04 & x06 & x09 & (x05 ? ~x02 : x08)))) | (x05 & ~x08 & ~x10 & ((~x02 & (x04 ? x06 : (~x06 & x09))) | (x02 & x04 & ~x06 & x09)))) : (~x04 & x05 & ((~x08 & (x02 ? (x06 ? (~x09 & x10) : x09) : (x06 ? (~x09 & ~x10) : (x09 & x10)))) | (x02 & ~x06 & x08 & x09 & x10)))) : (x05 ? ((x08 & ((x09 & ((~x03 & ((x02 & (x04 ? (x06 & x10) : ~x10)) | (x04 & ~x06 & x10))) | (~x02 & x03 & ~x04 & ~x06 & x10))) | (x03 & x04 & x06 & (x10 ? ~x09 : ~x02)))) | (x02 & ~x03 & x04 & ~x06 & ~x08 & x09 & ~x10)) : (x06 ? (x03 ? (x09 & ((x02 & x10 & (~x08 | (x04 & x08))) | (~x02 & x04 & x08 & ~x10))) : ((~x02 & ((~x04 & x08 & x09 & x10) | (x04 & ~x08 & ~x09 & ~x10))) | (x02 & ~x04 & ~x08 & ~x09 & ~x10))) : ((~x10 & ((x02 & ~x04 & (x03 ? (~x08 & x09) : (x08 & ~x09))) | (~x02 & x03 & x04 & ~x08 & x09))) | (~x08 & ~x09 & x10 & ~x02 & ~x03 & x04)))))) | (~x05 & x06 & ~x08 & ~x09 & ~x10 & x00 & x02 & x03 & x04))) | (~x02 & ((x04 & ((~x03 & ((x00 & ~x06 & x09 & x10 & (x01 ? (x05 & ~x08) : (~x05 & x08))) | (~x00 & x01 & x05 & x06 & ~x08 & ~x09 & ~x10))) | (~x06 & x08 & x09 & ~x10 & ~x00 & x01 & x03 & x05))) | (~x00 & x01 & x03 & ~x04 & x05 & x06 & x08 & ~x09 & ~x10)));
  assign z23 = (x04 & ((~x10 & ((~x07 & (x00 ? ((~x03 & ((x05 & ((x01 & ((~x06 & ~x08 & x09) | (x02 & x06 & x08 & ~x09))) | (x09 & ((~x02 & x06 & x08) | (~x01 & x02 & ~x08))))) | (x02 & ~x05 & x06 & x08 & ~x09))) | (~x02 & ((x03 & ((~x05 & ((x01 & x08 & (~x06 | (x06 & x09))) | (~x01 & x06 & ~x08 & ~x09))) | (~x01 & x05 & ~x06 & ~x09))) | (~x01 & ~x05 & ~x06 & ~x08 & x09)))) : (x02 ? (x01 ? (~x09 & ((~x03 & x06 & x08) | (~x06 & ~x08 & x03 & x05))) : (x05 & ((~x03 & x06 & x08) | (x03 & ~x06 & ~x08 & x09)))) : ((~x05 & ((~x06 & ((~x01 & x08 & (~x09 | (x03 & x09))) | (~x08 & x09 & x01 & x03))) | (~x01 & ~x03 & x06 & ~x08 & ~x09))) | (~x01 & x05 & x06 & ~x08 & x09))))) | (x07 & (x02 ? (x05 ? ((x00 & ~x09 & ((~x01 & ~x03 & x06) | (~x06 & x08 & x01 & x03))) | (~x00 & x01 & ~x03 & x06 & x08 & x09)) : ((x09 & (x00 ? (x03 & (x01 ? (~x06 & ~x08) : (x06 & x08))) : (~x03 & x08 & (x01 ^ x06)))) | (~x00 & ~x01 & ~x09 & (x03 ? (x06 & x08) : (~x06 & ~x08))))) : ((~x05 & ((~x08 & ((~x00 & x09 & ((~x03 & ~x06) | (~x01 & x03 & x06))) | (x00 & x01 & ~x03 & x06 & ~x09))) | (~x03 & x08 & ((~x01 & ~x06 & ~x09) | (x00 & (x01 ? (~x06 & ~x09) : (x06 & x09))))))) | (x05 & ~x06 & x08 & ~x00 & ~x01 & x03)))) | (x00 & ~x01 & ~x02 & ~x03 & x05 & ~x06 & x08 & ~x09))) | (x03 & (x08 ? (x10 & ((x01 & ((~x09 & ((x00 & ((x06 & (x02 ? (x05 ^ x07) : (~x05 & ~x07))) | (~x06 & x07 & ~x02 & x05))) | (~x00 & ~x02 & ~x05 & ~x06 & x07))) | (~x00 & ~x05 & ~x06 & x09 & (~x02 ^ x07)))) | (x00 & ~x01 & ((~x02 & ~x09 & (x05 ? (~x06 & ~x07) : (x06 & x07))) | (x02 & x05 & ~x06 & ~x07 & x09))))) : ((x10 & (x00 ? ((~x05 & ((x01 & ((~x02 & x06 & ~x07 & x09) | (x02 & ~x06 & x07 & ~x09))) | (~x01 & x02 & x06 & ~x07 & ~x09))) | (~x06 & x07 & x09 & ~x01 & ~x02 & x05)) : ((x01 & ((x09 & ((~x07 & (x02 ? (x05 ^ x06) : (x05 & x06))) | (~x02 & ~x05 & ~x06 & x07))) | (x05 & x06 & ~x09 & (~x07 | (x02 & x07))))) | (~x01 & x02 & x05 & ~x06 & x07 & x09)))) | (~x00 & ~x01 & x02 & ~x05 & x06 & ~x07 & x09)))) | (~x03 & (x00 ? ((x10 & ((~x09 & ((x05 & ((~x01 & ~x07 & ~x08 & (x02 ^ x06)) | (x07 & x08 & ((x02 & ~x06) | (x01 & ~x02 & x06))))) | (~x06 & x07 & x08 & ~x01 & ~x02 & ~x05))) | (x06 & x09 & ((x07 & ((x01 & (x02 ? (x05 & x08) : (~x05 & ~x08))) | (~x01 & x02 & ~x05 & ~x08))) | (x01 & ~x02 & ~x05 & ~x07 & x08))))) | (~x06 & ~x07 & x08 & x09 & ~x01 & ~x02 & ~x05)) : (x10 & ((x02 & ((x06 & (x01 ? (x05 & x08 & (x07 ^ x09)) : (~x08 & ((~x07 & x09) | (~x05 & x07 & ~x09))))) | (~x07 & x08 & ~x09 & x01 & x05 & ~x06))) | (x07 & ~x08 & ~x09 & x01 & ~x05 & x06))))))) | (~x04 & ((x10 & ((x01 & ((~x09 & (x00 ? ((x06 & ((~x02 & ~x05 & (x03 ? (~x07 & ~x08) : (x07 & x08))) | (x02 & x03 & x05 & x07 & x08))) | (x02 & ~x06 & x07 & (x03 ? (x05 & ~x08) : x08))) : (x02 ? ((~x06 & ~x07 & x03 & ~x05) | (x06 & x07 & ~x08 & ~x03 & x05)) : (x03 ? ((x06 & ~x07 & x08) | (x05 & x07 & ~x08)) : (x07 & (x05 ? (x06 & x08) : (~x06 & ~x08))))))) | (x09 & ((~x05 & x07 & ((~x00 & ((~x06 & x08 & ~x02 & x03) | (~x03 & x06 & ~x08))) | (x00 & ~x02 & ~x03 & ~x06 & x08))) | (x02 & x05 & ((x00 & ~x07 & ~x08 & (x03 ^ x06)) | (x06 & x08 & ~x00 & x03))))) | (x00 & x02 & ~x03 & x07 & ~x08 & ~x05 & x06))) | (x08 & ((~x01 & (x00 ? ((x02 & ~x05 & ((x03 & x07 & x09) | (~x03 & x06 & ~x07 & ~x09))) | (~x03 & x05 & x09 & ((x06 & x07) | (~x02 & ~x06 & ~x07)))) : ((x03 & ((x02 & x05 & ~x06 & ~x07 & x09) | (~x02 & ~x05 & x06 & x07 & ~x09))) | (~x03 & ((~x02 & ~x05 & ~x06 & ~x07 & x09) | (x02 & ((~x05 & x06 & x07 & x09) | (x05 & ~x06 & ~x07 & ~x09))))) | (~x02 & x05 & x06 & ~x07 & ~x09)))) | (x05 & ~x06 & ~x07 & ~x09 & ~x00 & ~x02 & x03))) | (~x01 & ~x08 & ((~x03 & ((~x05 & ((x07 & (x00 ? (~x09 & (x02 ^ x06)) : (~x06 & x09))) | (~x00 & x02 & x06 & ~x09))) | (x00 & ~x02 & x05 & x07 & x09))) | (x02 & x03 & x06 & x09 & (~x05 ^ x07)))))) | (~x10 & ((x02 & (x00 ? (x01 ? ((~x03 & x05 & ~x06 & x07 & x09) | (~x07 & ~x08 & ~x09 & x03 & ~x05 & x06)) : (~x05 & ((~x03 & ~x06 & ~x08 & (~x07 | (x07 & x09))) | (x08 & ~x09 & x03 & x07)))) : (x03 ? ((~x09 & ((~x01 & x05 & ~x08 & (x06 ^ ~x07)) | (~x07 & x08 & ~x05 & x06))) | (x07 & x08 & x09 & x01 & ~x05 & ~x06)) : (~x07 & ~x08 & ((~x01 & x05 & x06 & x09) | (x01 & (x05 ? x09 : (x06 & ~x09)))))))) | (~x08 & ((x07 & ((~x02 & ((x09 & ((x03 & (x00 ? ((x05 & ~x06) | (~x01 & ~x05 & x06)) : (~x01 & ~x05))) | (~x05 & ~x06 & ~x01 & ~x03))) | (~x00 & x01 & ~x03 & x05 & x06 & ~x09))) | (~x05 & x06 & ~x09 & ~x00 & x01 & x03))) | (~x02 & ~x07 & ((~x01 & ((x00 & ~x09 & (x03 ? (~x05 & ~x06) : (x05 & x06))) | (~x00 & ~x03 & ~x05 & x06 & x09))) | (x05 & ~x06 & ~x09 & x01 & x03))))) | (~x01 & ((~x02 & ((~x05 & ((~x06 & x08 & x09 & (x00 ? (x03 ^ x07) : (x03 & x07))) | (~x00 & x03 & x06 & ~x07 & ~x09))) | (~x07 & x08 & ~x09 & ~x03 & x05 & ~x06))) | (~x00 & ~x03 & ~x05 & x06 & x07 & x08 & x09))) | (~x00 & x01 & ~x02 & x03 & ~x07 & x08 & x05 & ~x06))) | (~x00 & x01 & x06 & x08 & ~x09 & ((~x05 & x07 & ~x02 & ~x03) | (x02 & x03 & x05 & ~x07))))) | (x00 & x10 & ((x01 & ~x02 & x06 & x08 & ((~x03 & ~x05 & ~x07 & ~x09) | (x03 & x05 & x07 & x09))) | (~x01 & x02 & x03 & ~x05 & ~x06 & ~x07 & ~x08 & x09)));
  assign z24 = (~x02 & ((~x00 & ((~x05 & ((x04 & (x01 ? ((x06 & ((x07 & ((~x03 & ~x10 & (x08 ^ ~x09)) | (x09 & x10 & x03 & ~x08))) | (x03 & ~x07 & x08 & (~x09 ^ x10)))) | (x03 & ~x06 & x07 & ~x08 & x09)) : ((~x07 & ((x03 & ((~x06 & x08 & x09 & ~x10) | (x06 & ~x08 & ~x09 & x10))) | (~x03 & ~x06 & ~x08 & ~x09 & ~x10))) | (~x06 & x07 & ~x09 & ((x08 & ~x10) | (~x03 & ~x08 & x10)))))) | (~x04 & (x03 ? (~x08 & ((~x06 & ~x07 & x09 & x10) | (x01 & ~x10 & (x06 ? (x07 & ~x09) : ~x07)))) : ((~x06 & ((x01 & ~x10 & ((~x08 & x09) | (~x07 & x08 & ~x09))) | (~x08 & x09 & x10 & ~x01 & x07))) | (~x01 & x06 & ((x07 & ~x08 & ~x09 & ~x10) | (~x07 & x08 & x09 & x10)))))) | (x07 & x08 & x09 & x10 & x01 & x03 & ~x06))) | (x05 & (x09 ? ((~x06 & ((x08 & x10 & ((~x01 & (x03 ? (~x04 & ~x07) : x07)) | (x01 & x03 & x04 & ~x07))) | (x01 & x04 & ~x10 & (x03 ? ~x07 : (x07 & ~x08))))) | (x03 & ((x10 & ((x01 & ~x04 & ((~x07 & ~x08) | (x06 & x07 & x08))) | (~x01 & x04 & x06 & ~x07 & ~x08))) | (~x07 & x08 & ~x10 & ~x01 & x04 & x06)))) : (x03 ? ((x04 & ((x07 & ((x06 & x08 & ~x10) | (~x01 & x10 & (~x06 | (x06 & x08))))) | (~x07 & ~x08 & ~x10 & ~x01 & ~x06))) | (x01 & ~x04 & ~x06 & ~x08 & x10)) : ((~x07 & ((x04 & x10 & (x01 ? x06 : (~x06 ^ x08))) | (x01 & ~x08 & ~x10 & (~x06 | (~x04 & x06))))) | (x01 & ~x06 & x07 & x08 & (~x04 ^ x10)))))) | (~x07 & x08 & ~x09 & x10 & ~x04 & x06 & x01 & x03))) | (x00 & ((x04 & ((x05 & (x06 ? (x03 ? ((~x01 & (x07 ? (~x08 & x09) : (x08 & ~x10))) | (~x08 & x09 & ~x10 & x01 & ~x07)) : (x07 & ((x01 & (x08 ? (~x09 & x10) : (x09 & ~x10))) | (x09 & x10 & ~x01 & ~x08)))) : ((x10 & ((~x07 & ((x01 & (x03 ? (x08 & ~x09) : (~x08 & x09))) | (~x01 & x03 & ~x08 & ~x09))) | (~x01 & x03 & x07 & x08 & x09))) | (x01 & ~x10 & ((~x07 & ~x08 & x09) | (~x03 & x07 & (x08 ^ ~x09))))))) | (~x05 & (x06 ? ((x09 & (x01 ? (~x10 & (x03 ? (x07 & ~x08) : (~x07 & x08))) : (x03 & x10 & (x07 ^ x08)))) | (~x01 & ~x03 & ~x09 & x10 & (x07 ^ x08))) : (x08 & ((~x07 & x09 & (x10 ? x03 : ~x01)) | (x07 & ~x10 & x01 & ~x03))))) | (x07 & x08 & ~x09 & x10 & ~x01 & ~x03 & ~x06))) | (~x04 & ((~x06 & (x10 ? ((x03 & ((~x05 & ~x07 & ~x08 & ~x09) | (x07 & (x01 ? (x08 & ~x09) : (x05 ? (x08 & ~x09) : (~x08 & x09)))))) | (x01 & ~x03 & ((~x05 & ~x07 & ~x08 & x09) | (x05 & x07 & x08 & ~x09)))) : ((~x01 & ((x03 & x05 & ((x08 & x09) | (x07 & ~x08 & ~x09))) | (~x03 & ~x05 & ~x07 & ~x08 & x09))) | (x01 & x03 & ~x05 & ~x07 & x08)))) | (x06 & ((x09 & ((x10 & ((x01 & ((~x03 & x07 & x08) | (~x07 & ~x08 & x03 & x05))) | (x07 & ~x08 & ~x03 & ~x05))) | (x07 & ~x08 & ~x10 & x03 & x05))) | (x08 & ~x09 & ~x10 & x03 & ~x05 & x07))) | (~x07 & ~x08 & ~x09 & ~x10 & x01 & ~x03 & ~x05))) | (~x07 & x08 & ~x09 & x10 & ~x05 & ~x06 & ~x01 & ~x03))) | (~x01 & ~x04 & ((~x03 & x08 & ((x05 & ~x06 & x07 & x09 & ~x10) | (~x05 & x06 & ~x07 & ~x09 & x10))) | (~x07 & ~x08 & x09 & x10 & x03 & ~x05 & x06))))) | (x02 & (x09 ? ((x01 & (x08 ? ((x05 & (x00 ? (x04 & x10 & (x03 ? (x06 ^ x07) : ~x06)) : (~x04 & ((~x06 & x07 & ~x10) | (~x07 & x10 & x03 & x06))))) | (x00 & ~x05 & ~x06 & ~x07 & (x03 ? (x04 & x10) : ~x04))) : (x10 ? (x03 ? ((~x00 & x04 & x05 & x06 & ~x07) | (x00 & ~x04 & x07 & (~x06 | (x05 & x06)))) : ((~x06 & ((~x00 & x05 & (~x04 ^ x07)) | (~x05 & ~x07 & x00 & x04))) | (~x00 & ~x04 & ~x05 & x06))) : ((x04 & (x00 ? (x03 & (x05 ? (x06 & x07) : (~x06 & ~x07))) : (~x03 & ~x05 & (x06 ^ x07)))) | (~x00 & x03 & ~x04 & ~x05 & x06 & x07))))) | (~x05 & ((~x01 & ((~x06 & ((x08 & (x00 ? ((~x04 & ~x07 & x10) | (x07 & ~x10 & x03 & x04)) : (x04 & x10 & (x03 ^ x07)))) | (x07 & ~x08 & x10 & x00 & ~x03 & ~x04))) | (x03 & ~x04 & x06 & ((x00 & ~x10 & (~x07 ^ x08)) | (~x08 & x10 & ~x00 & ~x07))))) | (x08 & ~x10 & x06 & x07 & x00 & ~x03 & x04))) | (~x01 & ((x05 & ((~x07 & ((x03 & ((x00 & ((x04 & x08 & ~x10) | (~x08 & x10 & ~x04 & ~x06))) | (~x00 & x04 & ~x06 & ~x08 & ~x10))) | (~x00 & ~x03 & x08 & (x04 ? (~x06 & x10) : (x06 & ~x10))))) | (~x00 & x06 & x07 & x10 & (x03 ? (~x04 & ~x08) : (x04 & x08))))) | (~x00 & x03 & ~x04 & x08 & ~x10 & ~x06 & ~x07)))) : ((x05 & (x01 ? (x03 ? ((~x07 & ((x00 & ((x08 & x10 & ~x04 & x06) | (~x08 & ~x10 & x04 & ~x06))) | (~x00 & ~x04 & x06 & ~x08 & ~x10))) | (~x00 & x07 & ((~x04 & x06 & ~x08 & x10) | (x08 & ~x10 & x04 & ~x06)))) : ((~x00 & ~x06 & ((~x04 & x08 & (x07 ^ ~x10)) | (x04 & x07 & ~x08 & ~x10))) | (~x07 & x08 & x10 & ~x04 & x06))) : (x08 ? ((~x06 & ((x00 & x04 & ~x10 & (~x07 | (~x03 & x07))) | (~x07 & x10 & ~x03 & ~x04))) | (x06 & ~x07 & x10 & x00 & x04)) : ((x04 & ((~x00 & ((~x03 & x06 & x10) | (x07 & ~x10 & x03 & ~x06))) | (x06 & ~x07 & ~x10 & x00 & x03))) | (~x03 & ~x04 & ((x06 & (x00 ? (~x07 | (x07 & x10)) : (x07 & ~x10))) | (x07 & x10 & ~x00 & ~x06))))))) | (~x05 & (x08 ? (x04 ? (x10 & ((~x00 & ((x06 & x07 & ~x01 & ~x03) | (x03 & ~x06 & ~x07))) | (x00 & ~x01 & x03 & ~x06 & x07))) : (x00 ? (~x03 & ((x06 & (x07 ? x01 : x10)) | (~x01 & ~x07 & ~x10))) : ((x07 & ((x10 & (x01 ? (x03 ^ x06) : (~x03 & ~x06))) | (~x01 & ~x03 & ~x10))) | (x06 & ~x07 & ~x10 & ~x01 & x03)))) : ((x10 & ((x03 & ((~x01 & ((x00 & x07 & (~x06 | (~x04 & x06))) | (~x00 & ~x04 & ~x06 & ~x07))) | (~x00 & x01 & x04 & x06 & x07))) | (x00 & ~x03 & x04 & ~x07 & (x01 ^ ~x06)))) | (~x06 & ~x07 & ~x10 & x01 & x03 & x04)))) | (~x00 & ~x01 & ~x04 & x06 & ((~x08 & ~x10 & ~x03 & ~x07) | (x08 & x10 & x03 & x07)))))) | (~x05 & ~x06 & ((~x00 & ~x07 & ~x08 & ((~x01 & ~x03 & ~x04 & ~x09 & x10) | (x01 & x03 & x04 & x09 & ~x10))) | (x00 & ~x01 & ~x03 & ~x04 & x07 & x08 & ~x09 & ~x10))) | (x00 & x01 & x03 & ~x04 & x05 & x06 & ~x10 & (x07 ? (x08 & x09) : (~x08 & ~x09)));
  assign z25 = (x10 & (x03 ? (x05 ? ((x02 & ((~x08 & (x06 ? ((x00 & x04 & (x01 ? (~x07 & ~x09) : (x07 & x09))) | (~x00 & x01 & ~x07 & x09)) : (x07 & ~x09 & (x01 ? ~x00 : ~x04)))) | (x01 & x08 & ((~x00 & ((~x04 & ~x06 & ~x07) | (x04 & x06 & x07 & x09))) | (x00 & x04 & ~x06 & ~x07 & ~x09))))) | (x04 & ((x01 & (x00 ? (~x02 & x07 & (x06 ? (x08 ^ ~x09) : (x08 & ~x09))) : ((~x06 & x07 & x08 & x09) | (~x02 & x06 & ~x07 & ~x08 & ~x09)))) | (~x02 & ~x06 & ~x07 & ~x09 & (x00 ? (~x01 & ~x08) : x08))))) : (x07 ? (((~x04 ^ x06) & ((x00 & x01 & x02 & x08 & x09) | (~x00 & ~x01 & ~x02 & ~x08 & ~x09))) | (x08 & ((~x01 & x02 & ~x04 & x06 & x09) | (~x00 & x01 & x04 & ~x06 & ~x09))) | (x02 & ((~x00 & x04 & ((~x01 & ~x06 & x09) | (~x08 & ~x09 & x01 & x06))) | (x00 & x01 & ~x04 & x06 & ~x08))) | (x00 & ~x02 & ~x04 & ~x08 & (x01 ? (~x09 | (~x06 & x09)) : (x06 & x09)))) : (x06 ? ((~x00 & ~x09 & ((x01 & ~x02 & x04 & x08) | (~x01 & x02 & ~x04 & ~x08))) | (x01 & x02 & x04 & ~x08 & x09)) : ((~x08 & ((x00 & ((~x01 & ~x02 & x04 & x09) | (x01 & x02 & ~x04 & ~x09))) | (~x00 & x01 & ~x02 & x04 & x09))) | (~x00 & ~x04 & x08 & (x01 ? (~x02 & x09) : ~x09)))))) : (x04 ? ((~x02 & ((~x01 & ((~x09 & ((~x05 & ~x06 & ~x07 & ~x08) | (x00 & x06 & (x05 ? ~x08 : (x07 & x08))))) | (~x00 & ~x06 & ~x07 & x09 & (x05 ^ x08)))) | (~x00 & ((x01 & ((x05 & ((~x06 & x07 & x08 & ~x09) | (x06 & ~x07 & ~x08 & x09))) | (~x05 & x06 & x07 & ~x08 & x09))) | (~x05 & x06 & ~x07 & ~x08 & x09))))) | (x05 & ((x09 & (x00 ? (~x07 & ((x06 & x08) | (x01 & x02 & ~x06 & ~x08))) : (x02 & x07 & ~x08 & (x01 ^ x06)))) | (~x00 & ~x01 & x02 & ~x06 & ~x07 & ~x08 & ~x09))) | (x07 & x08 & ((~x00 & x01 & x02 & x06 & x09) | (~x01 & ~x05 & ~x06 & ~x09)))) : (x02 ? ((x06 & ((x07 & ((x00 & ((~x01 & x05 & ~x09) | (x01 & ~x05 & ~x08 & x09))) | (~x00 & x01 & x05 & ~x08 & x09))) | (~x07 & x08 & ~x09 & ~x00 & x01 & ~x05))) | (~x01 & ~x06 & ((x00 & x09 & (x05 ? (x07 & x08) : (~x07 & ~x08))) | (x08 & ~x09 & x05 & ~x07)))) : (x08 ? (x05 ? (x06 & ((x00 & (x01 ? (x07 & x09) : (~x07 & ~x09))) | (~x00 & x01 & x07 & ~x09))) : ((~x01 & ((x00 & (x06 ? (x07 & x09) : (~x07 & ~x09))) | (~x00 & x06 & x07 & ~x09))) | (~x00 & x01 & ~x06 & x07 & x09))) : ((x01 & ~x09 & (x00 ? (x06 & (x05 ^ x07)) : (x05 & x07))) | (x06 & ~x07 & x09 & x00 & ~x01 & x05))))))) | (~x10 & (x06 ? (x04 ? (x01 ? (x00 ? ((~x08 & (x03 ? (~x09 & (x05 ? x02 : ~x07)) : ((~x05 & x07 & x09) | (~x02 & x05 & ~x07)))) | (~x02 & x03 & ~x07 & x08 & (x05 ^ ~x09))) : (~x09 & ((x02 & ~x03 & (x05 ? (~x07 & ~x08) : (x07 & x08))) | (~x02 & x03 & ~x05 & x07 & x08)))) : ((~x00 & ((~x02 & ~x03 & x05 & x07 & ~x08) | (x02 & x03 & ~x05 & ~x07 & x09))) | (x03 & ((x00 & ((x02 & ~x07 & ~x08 & (x05 ^ ~x09)) | (~x02 & x05 & x07 & x08 & x09))) | (~x02 & x05 & x07 & ~x08 & x09))) | (x02 & ~x03 & ~x08 & ((x05 & ~x07 & ~x09) | (x00 & ~x05 & x07 & x09))))) : (x00 ? (x02 ? (x01 ? ((~x03 & ~x05 & x07 & x08 & ~x09) | (x03 & x05 & ~x07 & ~x08 & x09)) : (~x03 & ~x05 & (x07 ? (x08 & x09) : (~x08 & ~x09)))) : (x07 & ~x09 & ((~x01 & ~x05 & x08) | (x03 & x05 & ~x08)))) : ((~x02 & ((x05 & (x01 ? (x03 & (x07 ? (~x08 & ~x09) : x08)) : (~x03 & (x07 ? (x08 & ~x09) : (~x08 & x09))))) | (x07 & x08 & x09 & ~x01 & x03 & ~x05))) | (~x01 & x02 & ~x03 & ~x05 & ~x07 & x08 & x09)))) : ((x07 & (x03 ? ((x02 & ((~x04 & ((x05 & ((~x00 & (x01 ? (x08 & ~x09) : (~x08 & x09))) | (x00 & x01 & x08 & x09))) | (~x00 & ~x01 & ~x05 & ~x08 & ~x09))) | (x00 & x08 & ((~x05 & x09) | (x01 & x04 & x05 & ~x09))))) | (~x02 & ((x00 & x08 & ((~x01 & ~x04 & x05 & x09) | (x04 & ~x05 & ~x09))) | (~x00 & x01 & ~x04 & ~x05 & ~x08 & x09))) | (~x05 & ~x08 & ~x09 & ~x00 & x01 & x04)) : ((~x02 & ((~x08 & ((~x00 & ((~x01 & ~x04 & ~x05) | (x01 & x04 & x05 & ~x09))) | (x00 & x01 & ~x04 & ~x05 & x09))) | (x05 & x08 & x09 & ~x00 & ~x01 & x04))) | (~x01 & x02 & ((x08 & ((x00 & ~x09 & (~x05 | (x04 & x05))) | (~x00 & ~x04 & ~x05 & x09))) | (~x00 & x04 & ~x08 & x09)))))) | (~x07 & ((~x04 & ((~x05 & (x00 ? (x03 & ((~x02 & ~x08 & ~x09) | (~x01 & x02 & x09))) : ((x01 & x08 & (x02 ? (~x03 & ~x09) : x09)) | (~x01 & x02 & ~x03 & ~x08 & x09)))) | (~x02 & x05 & ((x00 & x01 & (x03 ? (x08 & ~x09) : x09)) | (~x00 & ~x01 & x03 & x08 & x09))))) | (~x01 & x04 & ((~x08 & ((x03 & ~x09 & (x00 ? (~x02 | (x02 & x05)) : (x02 & ~x05))) | (~x00 & ~x02 & ~x03 & x05))) | (~x00 & x02 & ~x03 & ~x05 & x08 & x09))))) | (x00 & ~x01 & ~x02 & x03 & x08 & x09 & x04 & x05)))) | (x02 & ((~x03 & ~x09 & ((x00 & ~x05 & ((x06 & x07 & x08 & ~x01 & x04) | (~x06 & ~x07 & ~x08 & x01 & ~x04))) | (~x00 & ~x01 & ~x04 & x07 & ~x08 & x05 & ~x06))) | (~x00 & x03 & x09 & ((~x06 & x07 & x08 & ~x01 & x04 & x05) | (x01 & ~x04 & ~x05 & x06 & ~x07 & ~x08))))) | (x05 & ~x06 & ~x07 & ~x08 & ~x09 & ~x00 & ~x01 & ~x02 & x03 & ~x04);
  assign z26 = (x08 & (x03 ? ((~x10 & ((~x04 & (x01 ? (~x05 & ((x02 & x06 & ~x07 & ~x09) | (x00 & x07 & (x02 ? (~x06 & ~x09) : (x06 & x09))))) : (x00 ? ((~x02 & x05 & ~x06 & ~x07 & x09) | (x02 & ~x05 & x06 & x07 & ~x09)) : (x05 & ((~x02 & ~x06 & x07 & x09) | (x02 & x06 & ~x07 & ~x09)))))) | (x04 & ((~x05 & ((x01 & (x00 ? ((x02 & x07 & x09) | (~x02 & x06 & ~x07 & ~x09)) : (x06 & x07 & (x02 ^ x09)))) | (x00 & ~x01 & ~x07 & (x02 ? (x06 & x09) : (~x06 & ~x09))))) | (x00 & x05 & x07 & ((~x02 & ~x06 & x09) | (x01 & x02 & x06 & ~x09))))) | (x01 & x02 & ((x00 & ~x05 & x06 & ~x07 & x09) | (~x00 & x05 & ~x06 & x07 & ~x09))))) | (x10 & (x01 ? ((~x06 & ((x04 & ((x09 & (x00 ? (x02 & (~x05 ^ x07)) : (~x02 & ~x07))) | (~x00 & ~x02 & x05 & x07 & ~x09))) | (x02 & ((~x00 & ~x04 & ~x05 & ~x07 & x09) | (x00 & x05 & x07 & ~x09))))) | (x00 & x06 & ((x05 & ((x02 & ~x04 & (x07 ^ ~x09)) | (~x02 & x04 & x07 & ~x09))) | (x02 & ~x04 & ~x05 & ~x07 & x09)))) : ((x00 & ((x02 & x05 & ((x06 & x07 & ~x09) | (x04 & ~x06 & ~x07 & x09))) | (~x06 & x07 & ~x09 & ~x02 & x04 & ~x05))) | (x06 & ~x07 & ~x09 & x02 & x04 & ~x05)))) | (x05 & x06 & x07 & ~x09 & ~x02 & ~x04 & ~x00 & x01)) : (x00 ? (x06 ? ((x04 & (x01 ? ((x02 & ((x05 & ~x07 & ~x09) | (~x05 & x07 & x09 & x10))) | (~x02 & x05 & ~x07 & x09 & ~x10)) : (~x02 & ((~x05 & (x07 ? (~x09 & x10) : (x09 & ~x10))) | (x05 & x07 & x09 & ~x10))))) | (~x01 & ~x04 & ((x02 & ((x05 & x07 & x09 & ~x10) | (~x05 & ~x09 & (x07 ^ ~x10)))) | (~x02 & ~x05 & x07 & ~x09 & ~x10)))) : ((x04 & ((~x09 & ((x01 & ((x02 & ~x05 & x07) | (~x07 & ~x10 & ~x02 & x05))) | (~x01 & x02 & x05 & ~x07 & ~x10))) | (~x02 & x05 & x07 & x09 & x10))) | (x05 & x07 & x09 & ~x10 & x01 & x02 & ~x04))) : ((~x05 & (x01 ? (x02 ? (~x04 & ((x06 & x07 & ~x09 & x10) | (~x06 & ~x07 & x09 & ~x10))) : (x04 & x07 & (x06 ? ~x10 : (x09 & x10)))) : ((~x10 & ((x07 & ((~x04 & (x02 ? (x06 | (~x06 & x09)) : (~x06 & ~x09))) | (~x02 & x04 & x06 & x09))) | (~x02 & x04 & x06 & ~x07 & ~x09))) | (x02 & ~x04 & x09 & x10 & (x06 ^ ~x07))))) | (~x04 & ((x05 & ((~x07 & ((~x02 & (x01 ? (x06 & ~x09) : (x06 ? (x09 & ~x10) : (~x09 & x10)))) | (x01 & x02 & ~x10 & (~x06 ^ x09)))) | (x01 & ((~x02 & ~x06 & x09 & ~x10) | (x02 & x07 & x10 & (~x06 ^ x09)))))) | (x07 & x09 & x10 & ~x01 & ~x02 & ~x06))) | (x06 & ~x07 & x09 & x10 & x01 & x02 & x04 & x05))))) | (~x08 & ((~x02 & (x01 ? ((x00 & (x10 ? ((x06 & ((x03 & x07 & x09 & (x04 ^ x05)) | (~x03 & ~x04 & ~x05 & ~x07 & ~x09))) | (x03 & x04 & ~x06 & x07 & ~x09) | (~x03 & x05 & ~x07 & (x04 ? ~x09 : (~x06 & x09)))) : (x03 ? (~x04 & ~x07 & (x05 ? x06 : (~x06 & ~x09))) : (x04 & x07 & ~x09 & (x05 ^ ~x06))))) | (x03 & ((x07 & ((x04 & ((x05 & ~x06 & x09 & ~x10) | (~x05 & x06 & ~x09 & x10))) | (~x00 & ~x05 & ((x06 & ~x09 & ~x10) | (~x04 & x10 & (~x09 | (~x06 & x09))))))) | (~x00 & ~x04 & ~x07 & x09 & (x05 ? (x06 | (~x06 & x10)) : ~x10)))) | (x05 & x06 & x09 & x10 & ~x00 & ~x03 & ~x04)) : (x03 ? ((x06 & (x00 ? (~x09 & ((x04 & x07 & (~x05 | (x05 & x10))) | (~x07 & x10 & ~x04 & x05))) : ((x07 & x10 & ~x04 & x05) | (x04 & ~x05 & ~x07 & x09 & ~x10)))) | (~x07 & x09 & x10 & ~x00 & x04 & ~x06)) : ((~x06 & ((x09 & ((~x04 & ((x00 & x05 & (x07 ^ ~x10)) | (~x07 & ~x10 & ~x00 & ~x05))) | (~x00 & x04 & ~x05 & x07 & x10))) | (x05 & ~x09 & ((~x04 & ~x07 & ~x10) | (x07 & x10 & x00 & x04))))) | (x00 & ((~x04 & x05 & ~x07 & ~x09 & x10) | (x06 & ((x04 & ~x07 & ~x09 & (x05 ^ x10)) | (~x04 & ~x05 & x07 & x09 & ~x10))))))))) | (x02 & ((x09 & ((~x06 & ((~x10 & (x00 ? (~x03 & (x01 ? (~x04 & (x05 ^ x07)) : (~x07 & (~x05 | (x04 & x05))))) : (x03 & ((~x01 & (x04 ? (x05 & x07) : ~x05)) | (x04 & ~x05 & x07))))) | (~x03 & x04 & x10 & ((x00 & x05 & (x01 ^ x07)) | (~x05 & ~x07 & ~x00 & x01))))) | (~x03 & ((x06 & ((~x07 & ((x00 & ((x01 & ~x04 & ~x05) | (x05 & x10 & ~x01 & x04))) | (~x00 & ~x01 & ~x04 & ~x05 & x10))) | (~x00 & x01 & x07 & (x04 ? (x05 & ~x10) : (~x05 & x10))))) | (x05 & ~x07 & x10 & ~x00 & ~x01 & x04))) | (~x07 & x10 & ~x05 & x06 & x00 & x01 & x03 & x04))) | (~x09 & ((x04 & ((x05 & ((x00 & ~x06 & ((~x01 & ~x07 & x10) | (x07 & ~x10 & x01 & ~x03))) | (x06 & ~x07 & x10 & ~x00 & x01 & x03))) | (~x01 & ~x05 & ((~x00 & ((x03 & ~x07 & ~x10) | (x07 & x10 & ~x03 & x06))) | (~x06 & x07 & x10 & x00 & x03))))) | (x00 & x03 & ~x04 & ((~x01 & (x05 ? (x07 & (~x06 ^ ~x10)) : (~x07 & (~x06 ^ x10)))) | (~x06 & x07 & ~x10 & x01 & x05))))) | (x00 & x01 & x03 & x04 & x07 & ~x10 & ~x05 & x06))) | (~x09 & ((~x00 & ((~x01 & x03 & x04 & x05 & (x06 ? (~x07 & x10) : (x07 & ~x10))) | (x06 & x07 & ~x10 & x01 & ~x03 & ~x05))) | (~x05 & ~x06 & ~x07 & x10 & x00 & ~x01 & ~x03 & ~x04))))) | (~x00 & ((x01 & x05 & ~x06 & ((x07 & x09 & x10 & ~x02 & ~x03 & x04) | (~x07 & ~x09 & ~x10 & x02 & x03 & ~x04))) | (~x05 & x06 & x07 & ~x09 & x10 & ~x01 & x02 & x03 & ~x04)));
  assign z27 = (x01 & (x00 ? (x03 ? (x02 ? (x06 ? (x04 ? (x05 ? (x07 & (x08 ? (~x09 & ~x10) : x10)) : (~x07 & (x08 ? x10 : (x09 & ~x10)))) : (~x07 & ((~x05 & x08 & x09) | (x10 & (x05 ? (x08 ^ ~x09) : (~x08 & x09)))))) : ((~x04 & ~x10 & ((x08 & ~x09 & x05 & ~x07) | (~x05 & x07 & ~x08 & x09))) | (~x07 & x10 & ((x04 & x05 & ~x08) | (~x05 & x08 & x09))))) : (x09 ? ((~x10 & ((x05 & ((x07 & x08 & ~x04 & ~x06) | (~x07 & (x04 ? (x06 | (~x06 & x08)) : (~x06 & ~x08))))) | (x04 & ~x05 & x08 & (x06 ^ x07)))) | (~x06 & ((~x04 & x10 & (x05 ? (~x07 & x08) : (x07 & ~x08))) | (x07 & ~x08 & x04 & x05))) | (x07 & x08 & x10 & ~x04 & ~x05 & x06)) : ((x04 & x08 & ((~x05 & x07 & ~x10) | (~x07 & x10 & x05 & ~x06))) | (x07 & ~x08 & ~x10 & ~x04 & ~x05 & ~x06)))) : ((x10 & (x04 ? ((x08 & ((~x02 & ~x07 & (x05 ? (x06 & ~x09) : (~x06 & x09))) | (x07 & ((x02 & ~x06 & ~x09) | (x05 & x06 & x09))))) | (x02 & ~x05 & ~x08 & (x06 ? (~x09 | (x07 & x09)) : (~x07 & x09)))) : (x06 & (x02 ? ((~x05 & ~x07 & x08 & x09) | (x05 & x07 & ~x08 & ~x09)) : (x08 & (x05 ? (~x07 & x09) : (x07 & ~x09))))))) | (x09 & ((~x10 & ((x04 & (x02 ? ((~x07 & ~x08 & x05 & ~x06) | (x07 & x08 & ~x05 & x06)) : (~x06 & (x05 ? (x07 & x08) : (~x07 & ~x08))))) | (~x06 & x07 & ~x08 & ~x02 & ~x04 & x05))) | (x06 & ~x07 & x08 & ~x02 & ~x04 & ~x05))) | (~x06 & x07 & ~x09 & ~x10 & ((x02 & ~x05 & x08) | (~x02 & x04 & x05 & ~x08))))) : ((~x02 & (((x09 ^ x10) & ((x03 & ~x05 & ~x06 & (x04 ? (~x07 & ~x08) : x07)) | (x06 & ~x07 & ~x08 & ~x03 & ~x04 & x05))) | (x07 & (x05 ? (x03 ? ((x06 & x08 & ~x09 & ~x10) | (x04 & ~x06 & ~x08 & x09 & x10)) : (~x06 & ~x08 & ~x09 & (~x04 ^ x10))) : (x08 & ((~x03 & x04 & x06 & x10) | (~x04 & ~x06 & ~x09 & ~x10))))) | (~x07 & ((~x05 & ((~x03 & ((~x06 & ~x08 & x09 & x10) | (x08 & ~x10 & x04 & x06))) | (~x04 & x06 & x08 & ~x09 & x10))) | (x08 & x09 & ~x10 & ~x03 & x05 & ~x06))))) | (x02 & (x04 ? (x09 & x10 & ((~x07 & ((x03 & (x05 ? (~x06 & x08) : (x06 & ~x08))) | (x06 & x08 & ~x03 & ~x05))) | (x06 & x07 & x08 & ~x03 & x05))) : ((x07 & (x05 ? ((~x06 & ((~x03 & (x08 ? x10 : (x09 & ~x10))) | (~x09 & x10 & x03 & ~x08))) | (x03 & ~x10 & ((x08 & ~x09) | (x06 & ~x08 & x09)))) : (x09 & ((x03 & ~x08 & x10) | (x06 & ((~x08 & ~x10) | (~x03 & x08 & x10))))))) | (~x03 & ~x05 & ~x06 & ~x07 & x08 & x09)))) | (x07 & x08 & ~x09 & ~x10 & ~x05 & ~x06 & ~x03 & x04)))) | (~x01 & ((~x07 & (x08 ? (x00 ? ((~x10 & ((~x06 & ((~x02 & ~x03 & (x04 ? (~x05 & x09) : (x05 & ~x09))) | (x03 & ~x09 & ((x04 & x05) | (x02 & ~x04 & ~x05))))) | (x02 & x06 & ((x03 & x04 & x05) | (~x03 & ~x04 & ~x05 & x09))))) | (~x06 & x10 & ((~x02 & x03 & x04 & ~x05) | (x02 & ~x03 & ~x04 & x05 & ~x09)))) : ((~x05 & ((~x06 & ((~x02 & x03 & x04 & x09 & ~x10) | (x02 & ((~x03 & ~x04 & ~x10) | (x03 & x04 & x09 & x10))))) | (~x02 & ((~x03 & x04 & ((~x09 & x10) | (x06 & x09 & ~x10))) | (x03 & ~x04 & x06 & ~x09 & x10))))) | (x05 & x06 & ~x09 & x10 & ~x02 & ~x03 & x04))) : (x03 ? (x05 ? ((~x02 & ((x00 & ((x04 & x06 & x10) | (~x04 & ~x06 & ~x09 & ~x10))) | (~x00 & ~x04 & x06 & ~x09 & ~x10))) | (~x00 & x02 & x06 & (x04 ? (~x09 & x10) : (x09 & ~x10)))) : ((~x06 & ((x02 & ((x00 & x10 & (~x04 ^ x09)) | (~x00 & ~x04 & x09 & ~x10))) | (~x00 & ~x02 & ~x04 & x09 & x10))) | (~x02 & x04 & x06 & ((~x09 & x10) | (x00 & x09 & ~x10))))) : ((~x04 & (x09 ? ((~x00 & ~x10 & (x02 ? x06 : (~x05 & ~x06))) | (x02 & ~x05 & x06 & x10)) : ((x00 & ~x02 & (x05 ? (x06 & ~x10) : (~x06 & x10))) | (x02 & ((x05 & ~x06 & x10) | (~x00 & ~x05 & ~x10)))))) | (~x00 & x04 & ~x10 & ((x05 & x06 & ~x09) | (x02 & ~x05 & ~x06 & x09))))))) | (x07 & ((x08 & (x05 ? ((x06 & ((x10 & (x00 ? ((~x02 & ~x03 & ~x04) | (x02 & x03 & x04 & x09)) : (x03 & (x02 ? (~x04 & x09) : x04)))) | (~x02 & ~x03 & x04 & ~x09 & ~x10))) | (~x02 & ~x04 & ~x06 & x09 & (x00 ? x10 : ~x03))) : (x02 ? (x10 ? (x00 ? (x06 & (x03 ? (x04 & ~x09) : (~x04 & x09))) : (~x06 & (x03 ? (~x04 & x09) : (x04 & ~x09)))) : ((~x00 & (x03 ? (~x04 & ~x09) : (x04 & ~x06))) | (x04 & ~x06 & ~x09 & x00 & x03))) : ((~x09 & ((x00 & ~x03 & ~x04 & (~x06 ^ ~x10)) | (~x00 & x03 & x04 & x06 & ~x10))) | (x03 & x04 & ~x06 & x09 & x10))))) | (~x05 & ((~x08 & ((~x10 & ((x00 & ((x02 & ~x04 & x06 & x09) | (~x02 & ~x03 & x04 & ~x06 & ~x09))) | (x04 & x06 & ~x09 & ~x00 & ~x02 & ~x03))) | (~x00 & ((x04 & ((~x09 & x10 & (x02 ? (x03 | (~x03 & x06)) : ~x06)) | (~x02 & ~x03 & ~x06 & x09))) | (x02 & ~x03 & ~x04 & ~x06 & ~x09))))) | (~x04 & x06 & ~x09 & x10 & x00 & x02 & ~x03))) | (~x02 & x05 & ~x08 & ~x10 & ((~x00 & ((x03 & x09 & (~x04 ^ x06)) | (~x03 & x04 & ~x06 & ~x09))) | (x00 & x03 & ~x04 & x06 & ~x09))))) | (x00 & ~x02 & ~x03 & x04 & x05 & x06 & ~x08 & x09 & x10))) | (~x00 & x02 & x03 & x04 & ~x05 & ~x06 & ~x07 & x08 & ~x09 & x10);
  assign z28 = (~x05 & ((x07 & (x04 ? ((~x10 & (x00 ? ((x08 & ((~x01 & x03 & (x02 ? ~x09 : (~x06 & x09))) | (~x02 & ~x03 & x06 & x09))) | (x02 & ~x09 & (x01 ? (x03 & ~x08) : (~x03 & ~x06)))) : ((x08 & ((x06 & ~x09 & (x01 ? (x02 ^ ~x03) : (x02 & ~x03))) | (x01 & ~x02 & x03 & ~x06 & x09))) | (~x01 & ~x08 & (x02 ? (~x06 & x09) : (~x03 & ~x09)))))) | (x03 & ((x10 & ((~x00 & x09 & ((~x01 & x02 & x06 & x08) | (x01 & ~x02 & ~x06 & ~x08))) | (~x06 & x08 & ~x09 & x00 & x01 & x02))) | (~x00 & x01 & ~x02 & ~x06 & ~x08 & ~x09))) | (x00 & ~x01 & x02 & ~x03 & x08 & x10 & (~x06 ^ x09))) : ((x09 & (x02 ? (x01 ? (x10 & ((~x00 & ~x08 & (x03 ^ x06)) | (~x06 & x08 & x00 & x03))) : ((x08 & ((x00 & (x03 ? (x06 & ~x10) : (~x06 & x10))) | (x06 & ~x10 & ~x00 & ~x03))) | (~x08 & x10 & x00 & x06))) : ((x01 & ((~x08 & x10 & x03 & ~x06) | (x00 & ~x10 & (x03 ? (~x06 & x08) : (x06 & ~x08))))) | (~x00 & ~x01 & ~x06 & x08 & x10)))) | (~x09 & (x00 ? (x03 & ((x01 & x02 & x06 & (~x08 ^ ~x10)) | (~x01 & ~x02 & ~x06 & ~x08 & ~x10))) : ((~x06 & ((x01 & ((~x08 & x10 & ~x02 & ~x03) | (x02 & x03 & ~x10))) | (x08 & ~x10 & ((x02 & ~x03) | (~x01 & ~x02 & x03))))) | (~x01 & x02 & x03 & x06 & x08 & x10)))) | (~x00 & x01 & ~x02 & x08 & x10 & ~x03 & x06)))) | (~x02 & ((~x07 & (x04 ? (x00 ? ((~x06 & ((x09 & (x01 ? (x03 ? (x08 & x10) : (~x08 & ~x10)) : (~x08 & x10))) | (~x01 & x03 & ~x08 & ~x09 & ~x10))) | (x08 & ~x09 & ~x10 & x01 & x03 & x06)) : ((x06 & ((x01 & ~x10 & (x03 ? x09 : ~x08)) | (~x03 & x09 & x10 & (~x08 | (~x01 & x08))))) | (~x08 & x09 & x10 & ~x01 & x03 & ~x06))) : (x00 ? (x09 & ((x10 & ((x01 & ~x08 & (~x03 ^ x06)) | (x06 & x08 & ~x01 & ~x03))) | (x08 & ~x10 & x01 & ~x03))) : ((~x10 & ((~x03 & (x01 ? (x09 ? ~x08 : ~x06) : (x06 & ~x09))) | (~x01 & x03 & x06 & x08 & x09))) | (x08 & ~x09 & x10 & ~x01 & x03 & ~x06))))) | (x06 & ~x08 & ~x09 & x10 & x00 & ~x01 & x03 & ~x04))) | (x02 & ~x07 & (x03 ? ((x00 & x09 & ((~x04 & ((~x01 & (x06 ? (~x08 & ~x10) : (x08 & x10))) | (x08 & ~x10 & x01 & x06))) | (~x01 & x04 & x06 & ~x08 & x10))) | (~x00 & ~x01 & ~x04 & x06 & ~x08 & ~x09 & ~x10)) : (x01 ? ((x06 & ((x00 & ((x04 & x08 & ~x09) | (~x04 & ~x08 & x09 & x10))) | (x09 & ((~x04 & ~x08 & ~x10) | (~x00 & x04 & (x08 | (~x08 & x10))))))) | (x04 & ~x06 & ~x08 & ~x09 & ~x10)) : (~x06 & ((x04 & ((x00 & ~x08 & x10) | (~x00 & x08 & x09 & ~x10))) | (x00 & ~x04 & (x08 ? ~x09 : (x09 & x10)))))))))) | (x05 & (x02 ? (x04 ? (x08 ? (x01 ? (x09 ? (x00 ? (x06 & (x03 ? (x07 & ~x10) : ~x07)) : (~x06 & ~x10 & (x03 ^ ~x07))) : ((x00 & ~x03 & (x06 ? (~x07 & x10) : (x07 & ~x10))) | (x07 & x10 & x03 & x06))) : ((x03 & ((x00 & x10 & (x07 ? ~x06 : x09)) | (~x07 & ~x09 & ~x10 & ~x00 & ~x06))) | (x07 & ~x09 & x10 & x00 & ~x03 & x06))) : ((~x00 & ((x06 & (x01 ? ((x03 & ~x09 & ~x10) | (~x03 & x07 & x09 & x10)) : (x10 & (x09 ? (~x03 | (x03 & x07)) : ~x07)))) | (~x03 & ~x06 & ((x09 & x10 & x01 & ~x07) | (~x01 & ~x09 & ~x10))))) | (x00 & x07 & ((x09 & ~x10 & ~x01 & ~x06) | (x10 & ((x01 & (x03 ? ~x06 : (x06 & ~x09))) | (~x01 & ~x03 & ~x06 & x09))))) | (x01 & ~x03 & ~x06 & ~x07 & x09 & ~x10))) : (x03 ? ((x07 & ((~x08 & x09 & x10 & (x00 ? x01 : (x01 ^ ~x06))) | (x08 & ~x09 & ~x10 & ~x00 & ~x01 & ~x06))) | (~x00 & ~x01 & ~x07 & ((~x06 & ~x08 & ~x09 & ~x10) | (x06 & x08 & x09 & x10)))) : (x00 ? ((x07 & ((x01 & ~x08 & (x06 ? (x09 & ~x10) : (~x09 & x10))) | (x08 & ~x09 & x10 & ~x01 & ~x06))) | (~x08 & ~x09 & ~x10 & ~x01 & ~x06 & ~x07)) : ((x08 & ((x07 & ((x01 & (x06 ? (x09 & ~x10) : x10)) | (~x01 & x06 & x09 & x10))) | (~x01 & ~x06 & ~x07 & ~x09 & x10))) | (x01 & ~x08 & ((x06 & ~x07 & ~x09 & x10) | (~x06 & x07 & x09 & ~x10))))))) : ((x08 & (x01 ? (x04 ? ((~x07 & ((x00 & ~x10 & (x03 ? (~x06 & x09) : (x06 & ~x09))) | (~x00 & x03 & x06 & ~x09 & x10))) | (x07 & x09 & x10 & ~x00 & ~x03 & x06)) : (~x06 & ((~x00 & ~x03 & x07 & (~x10 | (x09 & x10))) | (~x09 & x10 & x03 & ~x07)))) : ((~x03 & ((~x06 & ((~x00 & ~x10 & (x04 ? (x07 & ~x09) : (~x07 & x09))) | (x09 & x10 & ~x04 & x07))) | (x07 & x09 & x10 & x00 & x04 & x06))) | (x00 & x03 & ~x04 & x06 & x10 & (x07 ^ x09))))) | (~x04 & ((x09 & ((~x03 & ((~x00 & ~x01 & ~x10 & (x06 ? ~x07 : (x07 & ~x08))) | (~x07 & ~x08 & x10 & x00 & x01 & x06))) | (x00 & x01 & ~x08 & ((~x06 & ~x07 & ~x10) | (x10 & ((~x06 & x07) | (x03 & (~x07 | (x06 & x07))))))))) | (x00 & ~x09 & x10 & ((x03 & (x01 ? (x06 ? ~x08 : x07) : (~x06 & ~x07))) | (~x01 & ~x03 & x06 & ~x07 & ~x08))))) | (x00 & x04 & ~x08 & (x06 ? ((~x07 & ((~x01 & x03 & x09 & ~x10) | (x01 & (x03 ? (~x09 & ~x10) : x10)))) | (~x01 & ~x03 & x07 & ~x09 & ~x10)) : ((~x01 & ~x03 & ~x07 & ~x09 & x10) | (x01 & x03 & x07 & x09 & ~x10))))))) | (~x01 & x04 & ~x06 & x09 & x10 & ((x00 & x03 & ~x08 & (x02 ^ x07)) | (~x00 & ~x02 & ~x03 & x07 & x08)));
  assign z29 = (~x02 & ((~x04 & ((x03 & ((~x10 & (x09 ? (x08 ? ((~x00 & ~x05 & (x01 ? (~x06 & ~x07) : x07)) | (x00 & ~x01 & x05 & ~x06 & ~x07)) : ((x01 & ((~x05 & ~x06 & ~x07) | (x00 & (x05 ? (~x06 & x07) : (x06 & ~x07))))) | (~x00 & ~x01 & x05 & x06 & x07))) : ((~x01 & ~x07 & (x00 ? (x05 & x06) : (~x06 & (x05 ^ x08)))) | (x06 & x07 & x08 & ~x00 & x01 & ~x05)))) | (x10 & (x06 ? ((~x00 & ((x01 & ((~x05 & x08 & x09) | (x05 & x07 & ~x08 & ~x09))) | (~x08 & ~x09 & ~x01 & x07))) | (x00 & ~x05 & x07 & x08 & x09)) : ((x07 & ((x05 & ((x00 & ((x08 & x09) | (x01 & ~x08 & ~x09))) | (~x00 & ~x01 & x08 & ~x09))) | (~x00 & x01 & ~x08 & x09))) | (x00 & ~x07 & x09 & (x01 ? (x05 & ~x08) : (~x05 & x08)))))) | (x00 & x01 & ~x05 & ~x06 & x07 & x08 & ~x09))) | (~x03 & (x07 ? ((~x06 & ((x05 & ((x01 & ((~x09 & x10 & ~x00 & ~x08) | (x09 & ~x10 & x00 & x08))) | (x00 & ~x01 & ~x09 & (~x10 | (~x08 & x10))))) | (x00 & ~x05 & x10 & ((~x08 & x09) | (~x01 & x08 & ~x09))))) | (x06 & x09 & x10 & x00 & ~x01 & x05)) : ((~x00 & (x01 ? (x09 & ((x08 & ~x10 & x05 & ~x06) | (x06 & ((~x08 & x10) | (~x05 & x08 & ~x10))))) : ((x09 & ((x05 & ~x10 & (~x06 ^ x08)) | (x08 & x10 & ~x05 & x06))) | (~x05 & ~x06 & ~x09 & (~x08 | (x08 & x10)))))) | (x09 & ((x05 & ((x00 & ((x01 & ~x08 & (~x06 ^ x10)) | (x08 & x10 & ~x01 & x06))) | (x08 & x10 & ~x01 & ~x06))) | (x00 & x01 & ~x05 & x06 & x08 & x10)))))) | (x07 & ~x08 & x09 & ~x10 & ~x05 & ~x06 & ~x00 & ~x01))) | (x04 & ((x05 & (x08 ? ((x01 & ((~x09 & ((x03 & x06 & (x00 ? (x07 & x10) : (~x07 & ~x10))) | (x00 & ~x03 & ~x06 & (~x10 | (~x07 & x10))))) | (x07 & ((~x00 & ((~x03 & ~x06 & ~x10) | (x03 & x06 & x09 & x10))) | (~x06 & x09 & x10 & x00 & x03))))) | (~x00 & ~x01 & x03 & ~x06 & ~x07 & x09 & x10)) : (x06 ? (x09 ? ((~x03 & ((x00 & (x01 ? x07 : (~x07 & x10))) | (~x00 & ~x01 & x07 & x10))) | (~x00 & x01 & x03 & (~x10 | (~x07 & x10)))) : ((~x00 & ~x01 & x07 & x10) | (x00 & ~x03 & ~x10 & (x01 ^ x07)))) : ((~x07 & ((x01 & ((x00 & ~x09 & (~x10 | (x03 & x10))) | (~x00 & ~x03 & x09 & x10))) | (~x00 & ~x01 & ~x03 & ~x09 & x10))) | (~x00 & ~x01 & ~x03 & x07 & x09 & ~x10))))) | (~x05 & (x07 ? ((~x00 & ((~x10 & (x01 ? (~x03 & (x06 ? (~x08 & ~x09) : x09)) : (x03 & x06 & (x08 ^ x09)))) | (~x06 & x10 & ((~x03 & x08 & ~x09) | (~x01 & x03 & x09))))) | (~x08 & ((x00 & x06 & ((~x03 & x09 & ~x10) | (~x01 & x03 & ~x09))) | (x01 & x03 & ~x06 & ~x09 & x10))) | (x00 & ~x01 & x06 & x08 & x09 & (~x10 | (~x03 & x10)))) : (~x08 & (x00 ? ((~x01 & ~x03 & ~x06 & ~x09 & ~x10) | (x06 & x09 & x10 & x01 & x03)) : (~x01 & x03 & ~x06 & (~x10 | (~x09 & x10))))))) | (x07 & x08 & ~x09 & ~x10 & x00 & x01 & x03 & x06))) | (x08 & ~x09 & ((~x00 & ~x03 & ~x05 & x07 & ~x10 & (x01 ^ x06)) | (x00 & ~x01 & x03 & x05 & x06 & ~x07 & x10))))) | (x02 & ((~x00 & (x10 ? (x07 ? (x01 ? ((~x08 & ((~x03 & ~x05 & ~x06 & (~x04 ^ x09)) | (x03 & x04 & x05 & x06 & ~x09))) | (~x06 & x08 & ~x09 & ~x03 & ~x04 & x05)) : (~x04 & ((x03 & ((~x06 & x08 & ~x09) | (x05 & ~x08 & x09))) | (~x03 & x05 & ~x06 & ~x09)))) : ((x01 & ((~x05 & (x03 ? (~x06 & (x04 ? (x08 & ~x09) : x09)) : (~x09 & (x04 ? ~x08 : (x06 & x08))))) | (x03 & x05 & x06 & (x04 ? (x08 & x09) : (~x08 & ~x09))))) | (~x01 & ((~x08 & ((~x05 & ((~x03 & ~x04 & x06 & ~x09) | (x03 & x04 & (~x06 ^ ~x09)))) | (~x03 & ~x04 & x05 & x09))) | (~x06 & x08 & x09 & ~x03 & x04 & x05))) | (~x03 & x04 & ~x05 & x06 & x08 & x09))) : (x08 ? (x03 ? ((x06 & ((~x01 & ((x04 & x05 & ~x07 & ~x09) | (~x04 & ~x05 & x07 & x09))) | (x01 & ~x04 & x05 & x07 & x09))) | (x01 & ((x04 & x05 & x07 & x09) | (~x04 & ~x06 & ~x09 & (~x05 ^ x07)))) | (~x04 & x05 & ~x06 & ~x07 & x09)) : ((~x04 & ((x01 & ((x05 & x06 & x07 & ~x09) | (~x05 & ~x06 & ~x07 & x09))) | (x07 & ~x09 & ~x01 & ~x06))) | (~x01 & x04 & ~x05 & x09 & (x06 ^ ~x07)))) : ((~x01 & ((x05 & ((x07 & ((~x03 & x04 & ~x06 & ~x09) | (x03 & (x04 ? x09 : (x06 & ~x09))))) | (~x03 & ~x04 & x06 & ~x07 & ~x09))) | (~x04 & ~x05 & x06 & ~x07 & ~x09))) | (~x04 & x09 & ((~x06 & x07 & x03 & ~x05) | (x01 & ~x03 & x05 & x06 & ~x07))))))) | (x00 & ((x05 & (x01 ? (x07 ? ((~x10 & ((x04 & ((x03 & (x06 ? (~x08 & x09) : (x08 & ~x09))) | (~x03 & ~x06 & x08 & x09))) | (~x03 & ~x04 & ~x06 & x08 & ~x09))) | (~x08 & ~x09 & x10 & x03 & ~x04 & x06)) : (x06 ? ((x08 & ~x10 & (x03 ? (~x04 ^ ~x09) : (x04 & x09))) | (~x08 & x10 & ~x03 & ~x04)) : ((~x03 & ~x04 & x08 & ~x09 & x10) | (x03 & x04 & ~x08 & x09 & ~x10)))) : ((~x03 & (x08 ? (x04 ? ((x06 & x07 & x09 & ~x10) | (~x06 & (x07 ? (~x09 & x10) : (x09 & ~x10)))) : ((~x06 & x07 & x09 & x10) | (x06 & ~x07 & ~x09 & ~x10))) : ((x06 & ~x07 & x09 & ~x10) | (~x06 & ((~x07 & ~x09 & x10) | (x04 & x07 & x09 & ~x10)))))) | (x03 & x04 & x06 & x07 & x08 & ~x10)))) | (~x05 & (x06 ? (x03 ? ((~x01 & x09 & ~x10 & (x04 ? (~x07 & x08) : (x07 & ~x08))) | (x08 & ~x09 & x10 & ~x04 & ~x07)) : ((~x07 & x08 & ~x09 & x01 & ~x04) | (x04 & ~x08 & ((x07 & ~x09 & ~x10) | (x01 & x10 & (x07 ^ x09)))))) : ((x07 & ((x10 & ((~x09 & (x01 ? (x08 & (x03 ^ ~x04)) : (~x03 & ~x04))) | (~x01 & ~x03 & x04 & ~x08 & x09))) | (~x01 & ~x03 & ~x04 & x08 & x09))) | (~x01 & x03 & x04 & ~x07 & x08 & x09 & x10)))) | (~x04 & ~x06 & x01 & x03 & x07 & x08 & x09 & ~x10))) | (~x06 & ~x07 & x08 & ~x09 & x10 & ~x04 & ~x05 & x01 & ~x03))) | (x00 & ~x07 & x08 & ~x10 & ((~x05 & ((x01 & ~x06 & ~x09 & (x03 ^ ~x04)) | (~x01 & x03 & ~x04 & x06 & x09))) | (x05 & ~x06 & ~x09 & ~x01 & x03 & x04)));
  assign z30 = (~x08 & ((~x09 & ((x07 & (x02 ? (x01 ? ((x04 & ((x00 & ~x10 & (x03 ? (x05 & x06) : (~x05 & ~x06))) | (~x00 & x03 & x05 & x06 & x10))) | (~x00 & ~x03 & ~x04 & x06 & (~x05 ^ x10))) : ((~x06 & x10 & ((~x03 & ~x04 & ~x05) | (~x00 & (x03 ? (~x04 & ~x05) : (x04 & x05))))) | (x05 & x06 & ~x10 & x00 & x03 & ~x04))) : (x00 ? (x01 ? ((~x03 & x04 & ~x05 & x06 & x10) | (x03 & ~x04 & ~x06 & ~x10)) : ((~x06 & (~x04 ^ x10) & (x03 ^ ~x05)) | (x03 & ~x04 & ~x05 & x06 & x10))) : ((~x01 & x06 & (~x03 ^ ~x04) & (~x05 ^ x10)) | (x05 & ~x06 & x10 & x01 & ~x03 & x04))))) | (~x07 & ((~x00 & (x05 ? ((x10 & ((x03 & ((x01 & (x02 ? (~x04 & x06) : (x04 & ~x06))) | (~x01 & x02 & x04 & x06))) | (~x02 & ~x03 & ~x04 & ~x06))) | (~x01 & ~x03 & ~x10 & (x02 ? (x04 & ~x06) : (~x04 & x06)))) : ((~x02 & ((x01 & x06 & (x03 ? x04 : (~x04 & x10))) | (~x01 & x03 & ~x04 & ~x06 & x10))) | (~x01 & x02 & x04 & ~x06 & x10)))) | (x05 & ((x00 & (x02 ? ((~x03 & x04 & x06 & ~x10) | (~x01 & ~x04 & x10 & (~x03 ^ x06))) : ((x01 & ((~x03 & ~x04 & ~x10) | (x03 & x04 & x06 & x10))) | (x04 & x06 & ~x01 & x03)))) | (~x06 & ~x10 & ((x01 & ~x02 & x03 & x04) | (~x01 & x02 & ~x03 & ~x04))))) | (~x03 & ~x05 & ~x06 & ~x10 & x00 & ~x01 & x02))) | (~x00 & x01 & x02 & x03 & x06 & x10 & x04 & ~x05))) | (x09 & (x10 ? (x01 ? ((~x05 & ((~x03 & ~x07 & ((x00 & (x02 ? x06 : (x04 & ~x06))) | (x04 & ~x06 & ~x00 & x02))) | (~x00 & ~x06 & x07 & (x02 ? (x03 & x04) : ~x04)))) | (x06 & ~x07 & x04 & x05 & ~x00 & ~x02 & ~x03)) : (x02 ? ((~x00 & ((x03 & x07 & ((x05 & ~x06) | (~x04 & ~x05 & x06))) | (~x03 & x04 & ~x05 & x06 & ~x07))) | (x05 & x06 & x07 & x00 & ~x03 & ~x04)) : ((x05 & ((~x06 & ((~x00 & ~x03 & ~x04 & ~x07) | (x00 & (x03 ? (~x04 & x07) : (x04 & ~x07))))) | (~x00 & ~x03 & ~x04 & x06 & x07))) | (~x05 & ~x06 & ~x07 & x00 & x03 & x04)))) : ((x02 & ((~x00 & ((x01 & ~x03 & ~x04 & x05 & x06) | (~x01 & x03 & x04 & ~x05 & ~x06 & ~x07))) | (x00 & ((x01 & ((x07 & ((x03 & (x04 ? (~x05 & ~x06) : (x05 & x06))) | (~x03 & x04 & ~x05 & x06))) | (~x03 & ~x04 & x06 & ~x07))) | (x05 & ~x07 & ((x03 & ~x04 & x06) | (x04 & ~x06 & ~x01 & ~x03))))) | (x01 & x03 & x04 & ~x05 & x06 & ~x07))) | (~x02 & ((x07 & (x03 ? ((~x00 & x01 & x04 & (x05 ^ ~x06)) | (x05 & x06 & ~x01 & ~x04)) : (x00 ? ((~x05 & x06 & ~x01 & x04) | (x05 & ~x06 & x01 & ~x04)) : (~x04 & x06 & (~x01 ^ x05))))) | (~x04 & ~x06 & ~x07 & (x00 ? (x01 ? (x03 & ~x05) : (~x03 & x05)) : (~x01 & ~x05))))) | (~x00 & x01 & ~x03 & ~x06 & x07 & x04 & ~x05)))) | (~x00 & x02 & ~x05 & x06 & ~x07 & ((~x04 & x10 & ~x01 & x03) | (x04 & ~x10 & x01 & ~x03))))) | (x08 & ((x04 & ((~x00 & ((~x03 & (x02 ? (x06 ? ((~x01 & ~x09 & (x05 ? (x07 & x10) : (~x07 & ~x10))) | (~x05 & ((x07 & x09 & ~x10) | (x01 & ~x07 & x10)))) : ((x07 & ((x01 & ~x09 & (~x10 | (x05 & x10))) | (~x01 & x05 & x09 & x10))) | (~x01 & ~x07 & (x05 ? (~x09 & x10) : (x09 & ~x10))))) : (x10 & ((~x05 & ((~x06 & ~x07 & ~x09) | (x01 & (x06 ? (~x07 & x09) : (x07 & ~x09))))) | (~x01 & x06 & (x09 ? x05 : ~x07)))))) | (x03 & ((~x02 & ((x05 & x06 & ~x07 & ~x09 & x10) | (x07 & x09 & ~x10 & ~x01 & ~x05 & ~x06))) | (x02 & ((x05 & x06 & x07 & x09 & ~x10) | (~x01 & x10 & ((x05 & ~x06 & ~x07 & x09) | (~x05 & x06 & x07 & ~x09))))) | (x07 & x09 & x10 & x01 & ~x05 & x06))) | (~x01 & x02 & ~x05 & ~x06 & ~x07 & ~x09 & ~x10))) | (x00 & (x03 ? ((~x02 & ((~x05 & ((x01 & ~x10 & (~x06 ^ x09)) | (~x01 & x06 & x07 & ~x09 & x10))) | (~x01 & x05 & x06 & x07 & x09 & ~x10))) | (x01 & x02 & x05 & ~x06 & x07 & ~x09 & ~x10)) : (x05 ? ((x01 & (x02 ? (x06 ? (x07 & ~x09) : (~x07 & x09)) : ((x06 & x07 & ~x09 & x10) | (~x06 & ~x10 & (x07 ^ ~x09))))) | (x07 & ~x09 & x10 & ~x01 & ~x02 & ~x06)) : ((x06 & ((~x01 & x07 & (x02 ? (x09 & x10) : (~x09 & ~x10))) | (x02 & ~x07 & ~x09 & x10))) | (~x01 & ~x02 & ~x06 & x09 & (x07 ^ x10)))))) | (x01 & x02 & x03 & ~x05 & x06 & x07 & ~x09 & ~x10))) | (~x04 & ((x02 & (x07 ? ((x01 & ((~x06 & ~x09 & x10 & x00 & ~x03 & x05) | (~x00 & x03 & ~x05 & x06 & x09 & ~x10))) | (~x01 & ((~x00 & ~x09 & (x03 ? (~x06 & ~x10) : (~x05 & x06))) | (x03 & ~x05 & ~x06 & x09 & x10))) | (x06 & ~x09 & ~x10 & ~x00 & x03 & x05)) : (x01 ? ((~x03 & ((~x00 & x09 & ((x06 & x10) | (~x05 & ~x06 & ~x10))) | (~x06 & ~x09 & ((x05 & x10) | (x00 & ~x05 & ~x10))))) | (x00 & x03 & x10 & (x05 ? (x06 & x09) : (~x06 & ~x09)))) : ((x06 & ((x00 & x05 & (x03 ? ~x10 : (x09 & x10))) | (~x00 & ~x03 & ~x05 & x09 & ~x10))) | (~x00 & ~x03 & ~x05 & ~x06 & x09 & x10))))) | (~x02 & ((x07 & ((~x09 & ((~x05 & ((~x00 & ((~x01 & ~x03 & x10) | (x06 & ~x10 & x01 & x03))) | (x00 & x01 & x03 & ~x06 & x10))) | (x00 & x05 & x10 & ((~x03 & ~x06) | (~x01 & x03 & x06))))) | (x01 & x05 & ~x06 & x09 & (x00 ? (~x03 & x10) : (x03 & ~x10))))) | (~x00 & ~x07 & ((x05 & ((x01 & x06 & (x03 ? (x09 & ~x10) : (~x09 & x10))) | (~x01 & x03 & ~x06 & x09 & x10))) | (x06 & ~x09 & ~x10 & ~x01 & x03 & ~x05))))) | (x06 & ~x07 & ~x09 & ~x10 & x00 & ~x01 & ~x03 & x05))) | (~x00 & ~x01 & ~x02 & ~x03 & x05 & x06 & x07 & ~x09 & ~x10))) | (x05 & ~x06 & x07 & x09 & ~x10 & x00 & ~x01 & x02 & x03 & x04);
  assign z31 = (x06 & (x02 ? ((x07 & ((x04 & ((x00 & ((x10 & ((x03 & ((~x01 & ~x09 & (x05 ^ x08)) | (x01 & ~x05 & x08 & x09))) | (x01 & ~x03 & ~x05 & (x08 ^ x09)))) | (x03 & x05 & ~x10 & (x01 ? (~x08 & x09) : (x08 & ~x09))))) | (~x00 & ((x01 & ~x10 & (x03 ? (x05 ? (x08 & ~x09) : x09) : (x08 & ~x09))) | (x08 & x09 & x10 & (x05 ? ~x03 : ~x01)))) | (~x08 & x09 & ~x10 & x01 & ~x03 & ~x05))) | (x03 & ((~x04 & ((~x08 & ((~x10 & ((x00 & ~x05 & (x01 ^ x09)) | (~x00 & x01 & x05 & x09))) | (~x00 & ~x01 & x05 & x09 & x10))) | (x08 & x09 & ~x10 & x00 & ~x01 & x05))) | (~x00 & ~x01 & x05 & ~x08 & ~x09 & x10))) | (~x04 & ~x05 & x08 & x09 & ~x10 & (x01 ? ~x00 : ~x03)))) | (x08 & (x04 ? (~x07 & ((x09 & ((~x00 & ((x01 & ~x05 & x10) | (~x01 & x03 & x05 & ~x10))) | (x00 & ~x01 & x03 & ~x05 & ~x10))) | (~x01 & ~x03 & x05 & ~x09 & ~x10))) : (x00 ? ((~x07 & ((x03 & ((x01 & x05 & (x09 ^ x10)) | (~x01 & ~x05 & ~x09 & x10))) | (~x01 & ~x03 & ~x05 & x09 & x10))) | (x01 & ~x03 & ~x05 & ~x09 & ~x10)) : (~x07 & x10 & ((x01 & x03 & (x05 ^ ~x09)) | (~x01 & ~x03 & x05 & ~x09)))))) | (~x08 & ((x03 & (x00 ? ((~x01 & ~x04 & x05 & x09 & x10) | (x04 & ~x05 & ~x07 & ~x09 & ~x10)) : (x05 & ~x07 & x09 & ~x10 & (~x01 ^ x04)))) | (~x07 & ((~x00 & ~x09 & ((x01 & x05 & x10) | (~x01 & ~x03 & x04 & ~x05 & ~x10))) | (x01 & ~x03 & ~x04 & x05 & x09 & x10)))))) : ((~x03 & ((x07 & (x00 ? (x09 ? ((~x01 & x04 & x05 & x08 & ~x10) | (x01 & x10 & (x04 ? (x05 & ~x08) : (~x05 & x08)))) : ((x04 & ((x05 & x08 & ~x10) | (x01 & x10 & (~x05 ^ x08)))) | (~x01 & ~x04 & ~x08 & (x05 ^ x10)))) : (~x04 & ((x01 & ((~x05 & x08 & ~x09 & ~x10) | (x05 & ~x08 & x09 & x10))) | (x09 & ~x10 & (~x05 ^ x08)))))) | (~x07 & ((x04 & ((x05 & ((~x00 & (x01 ? (~x09 & ~x10) : (x08 & x10))) | (x00 & ~x01 & ~x08 & ~x09 & x10))) | (x00 & ~x05 & x09 & ~x10 & (~x01 ^ x08)))) | (x00 & ~x04 & ~x09 & x10 & (x01 ? ~x08 : (x05 & x08))))) | (~x00 & ~x04 & x05 & ~x09 & (x01 ? (x08 & ~x10) : (~x08 & x10))))) | (x03 & (x04 ? ((~x08 & ((x00 & x01 & ~x05 & ((x09 & x10) | (x07 & ~x09 & ~x10))) | (~x01 & x05 & ((~x07 & ~x09 & ~x10) | (~x00 & (x07 ? (x09 & ~x10) : (~x09 & x10))))))) | (x05 & ((x00 & ((x09 & x10 & ~x01 & ~x07) | (x08 & ~x09 & ~x10 & x01 & x07))) | (x08 & x09 & x10 & ~x00 & ~x01 & x07))) | (~x07 & x08 & ~x09 & ~x10 & ~x00 & x01 & ~x05)) : ((x05 & ((x08 & ((~x00 & x10 & (x07 ? x09 : x01)) | (x00 & x01 & x07 & x09 & ~x10))) | (~x00 & x01 & ~x07 & ~x10 & (~x09 | (~x08 & x09))))) | (~x08 & ~x09 & x10 & ~x00 & ~x05 & ~x07)))) | (~x07 & ~x08 & ~x09 & x10 & ~x00 & ~x01 & x04 & ~x05)))) | (~x06 & (x09 ? ((x05 & (x02 ? ((~x03 & ((~x04 & ((~x00 & ~x10 & (x01 ? (x07 & x08) : (~x07 & ~x08))) | (x07 & x08 & x00 & ~x01))) | (x00 & x04 & (x01 ? (x07 & x10) : (x08 & ~x10))))) | (x00 & x01 & x03 & ~x08 & ~x10 & ~x04 & ~x07)) : (x00 ? (~x01 & ((~x08 & (x03 ? (x04 ? (x07 & ~x10) : (~x07 & x10)) : (x04 ? (~x07 & x10) : x07))) | (x07 & x08 & x03 & ~x04))) : ((x01 & ((~x03 & x07 & (x04 ? (x08 & x10) : (~x08 & ~x10))) | (x03 & ~x04 & ~x07 & ~x08 & x10))) | (x03 & x04 & ~x10 & (x08 ? ~x07 : ~x01)))))) | (~x05 & (x01 ? (~x02 & ((~x04 & ((~x00 & ~x03 & x08 & (x07 ^ ~x10)) | (~x08 & x10 & x03 & x07))) | (~x07 & ~x08 & ~x10 & ~x00 & ~x03 & x04))) : ((x10 & ((x04 & (x00 ? ((~x07 & x08 & x02 & ~x03) | (x07 & ~x08 & ~x02 & x03)) : (~x08 & (x02 ? x03 : (~x03 & ~x07))))) | (~x04 & x07 & x08 & x00 & x02 & ~x03))) | (~x04 & ~x10 & ((~x00 & ~x02 & (x03 ? (~x07 & ~x08) : (x07 & x08))) | (x07 & ~x08 & x00 & x03)))))) | (~x00 & ~x01 & x02 & ~x03 & x04 & x07 & ~x08 & ~x10)) : ((x05 & ((~x03 & (x01 ? ((x07 & ((x02 & ((x00 & ~x10 & (x04 | (~x04 & x08))) | (x08 & x10 & ~x00 & ~x04))) | (~x00 & ~x02 & x04 & ~x08 & x10))) | (x00 & ~x02 & ~x07 & (x04 ? (~x08 & x10) : (x08 & ~x10)))) : (x02 ? (~x08 & ~x10 & (x04 ? ~x00 : ~x07)) : (x10 & ((x00 & ~x07 & (x04 ^ ~x08)) | (x07 & x08 & ~x00 & x04)))))) | (x03 & (x01 ? (x07 & (x02 ^ x08) & ((~x04 & ~x10) | (x00 & x04 & x10))) : (x00 ? (x02 & ((~x07 & x08 & ~x10) | (~x08 & x10 & ~x04 & x07))) : (~x02 & ((x04 & x07 & ~x08 & x10) | (x08 & ~x10 & ~x04 & ~x07)))))) | (~x00 & x01 & ~x02 & x08 & x10 & ~x04 & ~x07))) | (~x05 & ((~x07 & ((x10 & ((~x02 & ((~x04 & (x00 ? (x01 ? (x03 & ~x08) : (~x03 & x08)) : (~x01 & ~x03))) | (~x00 & x01 & ~x03 & x04 & ~x08))) | (~x00 & x02 & ~x03 & x04 & (~x01 ^ x08)))) | (x04 & ~x10 & ((~x00 & ~x08 & (x01 ? (x02 & ~x03) : (~x02 & x03))) | (x00 & x02 & x03 & x08))))) | (x04 & x07 & ((x01 & ((~x00 & ~x02 & (x03 ? (~x08 & x10) : (x08 & ~x10))) | (x00 & x02 & x03 & ~x08 & ~x10))) | (~x01 & ~x02 & ~x03 & x08 & ~x10))))) | (x00 & x01 & x02 & ~x03 & x04 & x07 & x08 & x10)))) | (x00 & x01 & x02 & ~x03 & x04 & ~x05 & ~x07 & ~x08 & x09 & ~x10);
  assign z32 = (~x02 & ((~x10 & ((x09 & ((x00 & ((x04 & ((x03 & x05 & ~x06 & x07 & ~x08) | (x08 & ((~x06 & ~x07 & ~x01 & ~x05) | (x06 & ((x03 & (x01 ? (~x05 ^ x07) : (x05 & ~x07))) | (~x05 & x07 & ~x01 & ~x03))))))) | (~x04 & ((x07 & ~x08 & ((x01 & (x03 ? (~x05 & x06) : x05)) | (x05 & x06 & ~x01 & ~x03))) | (x06 & ~x07 & x08 & ~x01 & ~x03 & ~x05))) | (x06 & ~x07 & ~x08 & x01 & x03 & ~x05))) | (~x00 & ((~x07 & ((~x01 & x03 & x04 & (x05 ? (x06 ^ x08) : (x06 & x08))) | (~x05 & ~x06 & ~x08 & x01 & ~x03 & ~x04))) | (x05 & ((~x08 & ((x01 & x04 & (x03 ? ~x06 : (x06 & x07))) | (~x01 & x03 & ~x04 & x06 & x07))) | (~x06 & x07 & x08 & x01 & ~x03 & ~x04))))) | (~x01 & ~x03 & ~x04 & x07 & x08 & x05 & ~x06))) | (~x09 & (x07 ? ((~x05 & ((~x06 & ((x01 & x08 & (x00 ? x04 : (~x03 | (x03 & x04)))) | (~x04 & ~x08 & ~x01 & ~x03))) | (x00 & ~x01 & ~x03 & ~x08 & (x04 | (~x04 & x06))))) | (x00 & x05 & ((~x06 & x08 & ~x03 & ~x04) | (~x01 & (x03 ? (x06 & (x04 ^ ~x08)) : (~x04 & ~x08)))))) : ((x06 & (x00 ? (x01 & ((~x05 & x08 & x03 & ~x04) | (~x03 & x04 & x05 & ~x08))) : (~x01 & ((x03 & x05 & (~x08 | (x04 & x08))) | (~x05 & x08 & ~x03 & ~x04))))) | (x00 & ~x01 & x04 & ~x06 & ((x05 & x08) | (x03 & ~x05 & ~x08)))))) | (~x07 & x08 & x05 & ~x06 & x00 & x01 & x03 & ~x04))) | (x10 & (x09 ? ((~x07 & (x06 ? (~x08 & ((~x04 & ~x05 & x00 & x03) | (~x00 & ((x03 & ~x04 & x05) | (x04 & ~x05 & x01 & ~x03))))) : ((~x03 & ((x00 & ~x05 & (x01 ? (~x04 & ~x08) : (x04 & x08))) | (~x00 & ~x01 & x04 & x05))) | (~x00 & x03 & x05 & (x01 ? (x04 & x08) : ~x08))))) | (~x01 & ~x05 & x07 & ((x00 & ((~x03 & (x04 ? (~x06 & ~x08) : (x06 & x08))) | (x03 & x04 & x06 & ~x08))) | (~x00 & ~x03 & x06 & ~x08)))) : ((~x04 & (x06 ? ((x07 & ((~x05 & (x00 ? (x01 & ~x08) : (x08 & (x01 ^ x03)))) | (x00 & ~x01 & x05 & (~x03 ^ x08)))) | (~x00 & x01 & ~x08 & (x03 ? x05 : (~x05 & ~x07)))) : ((~x03 & ((~x01 & ((~x07 & ~x08 & ~x00 & x05) | (x00 & x08 & (x05 ^ x07)))) | (x05 & x07 & ~x00 & x01))) | (x00 & x01 & ~x05 & ~x07 & ~x08)))) | (~x07 & ((~x05 & ((x06 & ((x00 & ((~x01 & ~x08) | (x01 & ~x03 & x04 & x08))) | (~x00 & x01 & x03 & x04 & x08))) | (x04 & ~x06 & ~x08 & ((~x00 & ~x01 & ~x03) | (x01 & x03))))) | (x04 & x05 & ~x08 & ((x01 & ~x03 & ~x06) | (~x00 & ~x01 & x03 & x06)))))))) | (~x00 & x01 & ~x03 & x04 & x05 & ~x06 & ~x07 & x08 & x09))) | (x04 & ((x02 & (x06 ? (x00 ? (x03 ? ((~x08 & ((x01 & ~x09 & ~x10 & (x05 | (~x05 & x07))) | (~x01 & ~x05 & ~x07 & x09 & x10))) | (x08 & ~x09 & x10 & ~x01 & x05 & x07)) : (~x07 & ((x09 & x10 & (x01 ? (~x05 ^ x08) : (x05 & ~x08))) | (~x01 & x05 & x08 & ~x09 & ~x10)))) : (x05 ? ((x07 & ((x01 & x10 & (x03 ? (~x08 & ~x09) : (x08 & x09))) | (~x01 & x03 & x08 & ~x09 & ~x10))) | (x08 & x09 & ~x10 & ~x01 & ~x03 & ~x07)) : ((~x10 & ((~x01 & ~x08 & (x03 ? (~x07 & x09) : (x07 & ~x09))) | (x01 & ~x03 & ~x07 & x08 & ~x09))) | (x01 & x08 & x09 & x10 & (x03 ^ ~x07))))) : (x07 ? ((x08 & ((x00 & ((x09 & ((~x01 & x03 & x05 & ~x10) | (x01 & (x10 ? x05 : ~x03)))) | (~x01 & ~x03 & x05 & ~x09 & x10))) | (x05 & ~x09 & ~x10 & ~x00 & x01 & x03))) | (~x00 & ~x05 & ~x08 & x10 & (x01 ? (~x03 ^ x09) : (~x03 & x09)))) : ((x00 & ~x08 & (x01 ? ((~x03 & ~x05 & ~x09 & x10) | (x03 & x05 & x09 & ~x10)) : (x05 & (x03 ? (~x09 & x10) : (x09 & ~x10))))) | (~x01 & x03 & x05 & x08 & x09 & x10))))) | (x00 & x03 & x06 & x10 & ((x01 & x05 & (x07 ? (x08 & ~x09) : (~x08 & x09))) | (~x01 & ~x05 & x07 & x08 & ~x09))) | (~x06 & ~x07 & ~x08 & x09 & ~x10 & ~x00 & ~x01 & ~x03 & x05))) | (x02 & ((~x04 & (x00 ? (x08 ? ((~x07 & ((~x06 & (x03 ? ((x01 & (x05 ? x10 : (~x09 & ~x10))) | (~x01 & x05 & ~x09 & ~x10)) : (~x05 & ((~x09 & ~x10) | (~x01 & x09 & x10))))) | (~x03 & ~x05 & x06 & ~x09 & (~x01 ^ x10)))) | (~x03 & x07 & (x01 ? ((~x05 & ~x06 & x09 & x10) | (x05 & x06 & ~x09 & ~x10)) : (x06 & x10 & (~x05 | (x05 & x09)))))) : ((x06 & ((x05 & ((~x03 & ~x07 & x09 & ~x10) | (~x01 & ~x09 & (x03 ? (~x07 & x10) : (x07 & ~x10))))) | (x03 & ~x05 & ~x09 & ((~x07 & x10) | (~x01 & x07 & ~x10))))) | (~x01 & x03 & x05 & ~x06 & x07 & ~x09 & ~x10))) : ((x05 & (x01 ? (~x03 & ((~x06 & ~x07 & ~x09 & ~x10) | ((x06 ? (~x07 & ~x10) : (x07 & x10)) & (x08 ^ x09)))) : (x03 & x06 & ~x08 & (x07 ? (~x10 | (x09 & x10)) : (x09 & ~x10))))) | (x01 & x03 & ~x05 & ((~x10 & ((~x06 & ~x07 & ~x08 & ~x09) | (x06 & x07 & (x08 ^ x09)))) | (~x06 & ~x07 & x08 & x09 & x10)))))) | (x00 & x01 & ~x03 & x05 & ~x06 & ~x07 & ~x08 & x09 & x10)));
  assign z33 = (~x00 & ((x08 & ((x04 & (((x03 ^ ~x07) & ((x01 & ~x06 & ((x02 & x05 & ~x09 & x10) | (~x02 & ~x05 & x09 & ~x10))) | (~x01 & x02 & x05 & x06 & x09 & ~x10))) | (~x01 & ((~x09 & ((~x06 & ((~x03 & ~x10 & (x02 ? (x05 ^ x07) : (x05 & x07))) | (~x02 & x03 & ~x05 & ~x07 & x10))) | (x02 & ~x03 & x06 & x07 & (x05 ^ x10)))) | (x05 & x09 & x10 & ((~x03 & ~x06 & x07) | (x02 & x03 & x06 & ~x07))))) | (x01 & x02 & x03 & x09 & ((~x05 & x10 & (x06 ^ x07)) | (~x10 & ((x06 & ~x07) | (x05 & ~x06 & x07))))))) | (~x04 & (x01 ? (x06 ? ((~x03 & ((~x07 & ((x02 & ((x09 & ~x10) | (~x05 & ~x09 & x10))) | (x09 & x10 & ~x02 & x05))) | (~x02 & x05 & x07 & ~x09 & x10))) | (x02 & ~x05 & x07 & ~x10 & (~x09 | (x03 & x09)))) : ((x02 & x07 & ~x09 & (x03 ? (x05 & ~x10) : (~x05 & x10))) | (~x02 & x03 & ~x05 & x09 & ~x10))) : (x05 ? ((~x09 & ((x03 & ((x02 & (x06 ? (x07 & x10) : ~x07)) | (x07 & ~x10 & ~x02 & x06))) | (x07 & x10 & ~x02 & ~x03))) | (~x07 & x09 & ~x10 & ~x02 & ~x03 & ~x06)) : (x06 & (x03 ? (x09 & (x02 ? (~x07 & ~x10) : (x07 ^ x10))) : ((~x07 & x09 & ~x10) | (~x02 & x07 & x10))))))) | (x06 & ((~x09 & ((x01 & x07 & ((x02 & x03 & ~x05 & x10) | (~x02 & ~x03 & x05 & ~x10))) | (~x01 & ~x02 & ~x03 & x05 & ~x07 & ~x10))) | (~x01 & ~x02 & x03 & x09 & ~x10 & x05 & ~x07))))) | (~x08 & (x07 ? ((x06 & (x03 ? ((~x04 & ((x01 & ~x09 & ~x10 & (x02 ^ ~x05)) | (~x01 & ~x02 & x05 & x09 & x10))) | (~x01 & x10 & ((~x02 & ~x05 & x09) | (x02 & x04 & x05 & ~x09)))) : (x04 & ((x05 & ((x01 & x10 & (x02 | (~x02 & x09))) | (~x01 & x02 & x09 & ~x10))) | (~x01 & x02 & ~x05 & ~x09))))) | (x03 & ((x01 & x09 & x10 & ((x02 & ~x04 & ~x05) | (~x02 & x04 & x05 & ~x06))) | (~x05 & ~x09 & ~x10 & ~x01 & x02 & x04)))) : ((x01 & ((x04 & ((~x06 & (x02 ? ((x03 & x05 & x10) | (~x03 & ~x05 & ~x09 & ~x10)) : ((~x05 & x09 & ~x10) | (~x03 & (x05 ? (x09 & ~x10) : (~x09 & x10)))))) | (~x02 & x03 & x05 & x06 & x09 & x10))) | (~x02 & ~x04 & ((x03 & ((x05 & x09 & x10) | (~x05 & ~x06 & ~x09 & ~x10))) | (~x03 & ~x05 & x06 & x09 & ~x10))))) | (x05 & x06 & x09 & x10 & x02 & ~x03 & x04) | (~x01 & ((x09 & ((x03 & ~x10 & ((x05 & x06 & x02 & ~x04) | (~x05 & ~x06 & ~x02 & x04))) | (~x02 & ~x03 & x05 & x10 & (x04 ^ x06)))) | (x06 & ~x09 & ((x02 & ~x03 & ((x05 & x10) | (~x04 & ~x05 & ~x10))) | (~x02 & ~x04 & ~x05 & x10)))))))) | (~x01 & x03 & x04 & ~x07 & x10 & ((x02 & ~x05 & x06 & x09) | (~x02 & x05 & ~x06 & ~x09))))) | (x00 & ((~x03 & ((~x08 & (x01 ? (x02 ? (x06 & ((x04 & ((x05 & (x07 ? ~x09 : (x09 & x10))) | (~x05 & x07 & ~x09 & x10))) | (~x04 & ~x05 & ~x07 & ~x09 & x10))) : (x04 ? (x09 & ((x07 & ~x10 & ~x05 & x06) | (~x07 & x10 & x05 & ~x06))) : (~x06 & ~x07 & ~x09 & (~x05 ^ x10)))) : ((x10 & ((~x02 & ((~x04 & ~x05 & ~x06 & ~x07 & x09) | (x04 & x05 & x06 & x07 & ~x09))) | (x02 & ((x04 & ((~x05 & x07 & x09) | (x05 & ~x06 & ~x07 & ~x09))) | (~x04 & x05 & x06 & x07 & ~x09))) | (~x04 & ~x05 & ~x06 & x07 & ~x09))) | (x05 & ~x10 & ((~x02 & ~x06 & (x04 ? (x07 & ~x09) : (~x07 & x09))) | (x02 & x04 & x06 & ~x07 & ~x09)))))) | (x08 & (x07 ? (x09 ? ((~x04 & ((x05 & x10 & (x01 ? (~x02 | (x02 & x06)) : x06)) | (~x01 & x02 & ~x06 & ~x10))) | (~x01 & x04 & x06 & (x02 ? (~x05 & ~x10) : (x05 & x10)))) : (x10 & ((x01 & ~x06 & (x02 ? (x04 & ~x05) : x05)) | (~x01 & ~x02 & x04 & ~x05 & x06)))) : (x01 ? (x02 & x06 & ((x04 & ~x05 & ~x09) | (~x04 & x05 & x09 & ~x10))) : (~x06 & x09 & x10 & ((x04 & ~x05) | (~x02 & ~x04 & x05)))))) | (x06 & ~x07 & ~x09 & x10 & ~x01 & ~x02 & ~x04 & x05))) | (x03 & ((x05 & (x07 ? ((~x04 & ((x09 & ((x02 & ((~x06 & x08 & x10) | (~x08 & (x01 ? (~x06 ^ x10) : (x06 & ~x10))))) | (x08 & x10 & ~x02 & x06))) | (~x01 & ~x02 & ~x06 & ~x09 & ~x10))) | (~x01 & x04 & ((x02 & x06 & ~x08 & ~x09) | (~x02 & ~x06 & x08 & x09 & x10)))) : (x01 ? ((~x10 & ((x09 & ((x02 & (x04 ? (~x06 & x08) : (x06 & ~x08))) | (~x06 & ~x08 & ~x02 & ~x04))) | (~x02 & x04 & x06 & ~x08 & ~x09))) | (x02 & ~x04 & ~x06 & x09 & x10)) : (~x02 & ~x04 & x10 & ((~x06 & x08 & ~x09) | (~x08 & (~x09 | (x06 & x09)))))))) | (~x05 & (x08 ? (x01 ? ((x04 & x10 & (x02 ? (~x06 & ~x09) : (x07 & x09))) | (~x02 & ~x04 & ~x09 & ~x10 & (x06 ^ x07))) : ((x04 & x06 & ((x02 & ~x07 & ~x09 & x10) | (~x02 & x07 & x09 & ~x10))) | (x02 & ~x04 & ~x06 & ~x07 & (x09 ^ x10)))) : ((~x04 & ((x01 & ~x06 & ~x09 & x10 & (~x02 ^ x07)) | (~x01 & ~x02 & x06 & x09 & ~x10))) | (~x01 & x02 & x04 & ~x06 & x07 & ~x09 & x10)))) | (x07 & x08 & ~x09 & ~x10 & x01 & x02 & x04 & x06))) | (x04 & ~x06 & ((x02 & x05 & ((x08 & x09 & x10 & ~x01 & ~x07) | (x01 & x07 & ~x08 & ~x09 & ~x10))) | (~x01 & ~x02 & ~x05 & x08 & (x07 ? (x09 & x10) : (~x09 & ~x10))))))) | (~x03 & ~x08 & ((x06 & ~x07 & ((~x01 & x04 & ~x05 & (x02 ? (x09 & ~x10) : (~x09 & x10))) | (x05 & ~x09 & ~x10 & x01 & x02 & ~x04))) | (~x06 & x07 & ~x09 & x10 & ~x01 & ~x02 & ~x04 & x05)));
  assign z34 = (x04 & ((x00 & ((~x09 & (x10 ? ((~x07 & (x02 ? (x01 ? ((x03 & ~x05 & (~x06 | (x06 & x08))) | (~x06 & x08 & ~x03 & x05)) : ((~x03 & x05 & ~x08) | (~x06 & x08 & x03 & ~x05))) : ((~x01 & x03 & (x05 ? (~x06 & x08) : (x06 & ~x08))) | (x06 & ~x08 & x01 & x05)))) | (~x03 & x07 & (x01 ? (~x08 & (x02 ? x05 : (~x05 & ~x06))) : (x08 & (x02 ? (x05 & x06) : (~x05 & ~x06)))))) : (x01 ? (~x05 & ((~x02 & ((~x03 & ~x06 & x07) | (~x07 & ~x08 & x03 & x06))) | (x02 & ~x03 & ~x06 & ~x07 & x08))) : ((x02 & ((~x06 & ((x03 & (x05 ? x07 : (~x07 & ~x08))) | (x07 & x08 & ~x03 & ~x05))) | (~x03 & ~x05 & x06 & (x07 ^ x08)))) | (~x02 & ~x03 & x05 & x07 & x08))))) | (x03 & ((x09 & ((x06 & ((~x01 & ((x02 & ~x05 & x07 & ~x08 & x10) | (~x07 & x08 & ~x10 & ~x02 & x05))) | (x01 & x02 & ~x05 & ~x07 & ~x08 & x10))) | (x01 & ~x06 & ((~x07 & ((x05 & ~x08 & ~x10) | (x02 & x08 & (~x05 ^ x10)))) | (x07 & ~x08 & x10 & ~x02 & x05))))) | (x02 & x05 & x06 & x07 & (x01 ? (~x08 & x10) : (x08 & ~x10))))) | (x09 & ((~x03 & ~x10 & ((~x06 & ((~x07 & ((x01 & ((~x05 & ~x08) | (x02 & x05 & x08))) | (~x01 & x02 & x05 & ~x08))) | (x01 & ~x02 & ~x05 & x07 & x08))) | (x06 & ~x07 & ~x08 & x01 & ~x02 & x05))) | (~x08 & x10 & ~x06 & ~x07 & x01 & ~x02 & x05))))) | (~x00 & (x03 ? ((~x01 & (x07 ? (~x10 & ((x02 & ~x05 & x06 & x08 & ~x09) | (~x02 & (x05 ? (~x08 & x09) : (~x06 & ~x09))))) : ((x05 & ((~x06 & x08 & ~x10) | (x02 & x09 & (x06 ? (~x08 & ~x10) : (x08 & x10))))) | (~x02 & ~x05 & ((x06 & x08 & ~x09 & ~x10) | (~x08 & ((~x09 & ~x10) | (~x06 & x09 & x10)))))))) | (x01 & (x05 ? ((x07 & ~x09 & ((x06 & x08 & ~x10) | (~x08 & x10 & ~x02 & ~x06))) | (~x02 & x06 & ~x07 & x09 & (~x08 ^ ~x10))) : ((~x06 & ((~x07 & x08 & ~x09 & ~x10) | (~x02 & x07 & ~x08 & x09 & x10))) | (x02 & x06 & x07 & ~x09 & x10)))) | (x07 & x08 & ~x09 & ~x10 & ~x02 & x05 & ~x06)) : (x08 ? (x05 ? ((~x06 & ((~x09 & ((x01 & x02 & (x07 ^ ~x10)) | (~x01 & ~x02 & x07 & x10))) | (~x02 & ~x07 & x09 & ~x10))) | (~x01 & x06 & ~x10 & (x02 ? (x07 & ~x09) : x09))) : (~x09 & ((~x01 & ((~x07 & x10 & ~x02 & x06) | (x02 & ~x06 & (x07 ^ ~x10)))) | (x01 & ~x02 & x06 & ~x07 & ~x10)))) : ((x01 & x07 & ((x05 & ((~x06 & ~x09) | (x02 & x06 & x09 & x10))) | (x02 & x09 & ((~x06 & x10) | (~x05 & x06 & ~x10))))) | (~x07 & x09 & x10 & ~x01 & ~x05 & ~x06))))) | (x06 & x07 & x08 & ((~x01 & ~x02 & ~x05 & x10 & (x03 ^ x09)) | (x05 & x09 & ~x10 & x01 & x02 & x03))))) | (~x04 & ((x03 & ((~x10 & (x05 ? (x00 ? (x06 & ((~x08 & ((x07 & (x01 ? (x02 | (~x02 & x09)) : (x02 & x09))) | (~x01 & x02 & ~x07 & ~x09))) | (x01 & ~x02 & ~x07 & x08 & ~x09))) : ((~x01 & x08 & x09 & (x02 ? (~x06 & x07) : (x06 & ~x07))) | (x01 & ~x02 & ~x06 & ~x07 & ~x08))) : (x01 ? ((x00 & ((x02 & x06 & ~x07 & ~x09) | (~x02 & ~x06 & x07 & x08 & x09))) | (x07 & ~x08 & ~x09 & ~x00 & x02 & ~x06)) : ((~x07 & ((~x06 & ((x00 & (x08 ? x09 : ~x02)) | (x02 & ~x08 & x09))) | (~x00 & x06 & (x02 ? (x08 & ~x09) : ~x08)))) | (x00 & ~x02 & x06 & x07 & x08))))) | (x10 & ((~x09 & (x01 ? (~x05 & ((~x00 & ~x06 & ~x08 & (x02 ^ x07)) | (x00 & x02 & x06 & x07 & x08))) : ((x02 & x08 & ((x00 & ~x07 & (x05 ^ x06)) | (x06 & x07 & ~x00 & x05))) | (~x00 & ~x02 & ~x08 & (x05 ? x07 : (~x06 & ~x07)))))) | (~x08 & x09 & ((~x02 & ((~x00 & ((x01 & ~x07 & (x05 ^ x06)) | (x06 & x07 & ~x01 & x05))) | (x00 & ~x01 & ~x05 & ~x06 & x07))) | (~x00 & x01 & x02 & ~x06 & x07))))) | (x02 & ~x05 & x06 & x09 & ((~x07 & x08 & x00 & ~x01) | (x07 & ~x08 & ~x00 & x01))))) | (~x03 & (x06 ? (x05 ? ((x02 & (x00 ? (x10 & ((x01 & x07 & (x08 ^ ~x09)) | (x08 & ~x09 & ~x01 & ~x07))) : (~x10 & ((x07 & x08 & x09) | (x01 & ~x08 & ~x09))))) | (x00 & ~x09 & x10 & (x01 ? (~x07 & x08) : (~x02 & x07)))) : ((~x02 & ((x00 & x08 & x09 & (x01 ? (x07 & ~x10) : (~x07 & x10))) | (~x08 & ~x09 & x10 & ~x01 & x07))) | (x00 & ~x01 & x02 & ~x07 & ~x08 & x09 & x10))) : (x10 ? (x00 ? ((x01 & ~x08 & ((x05 & ~x07 & ~x09) | (x02 & ~x05 & x07 & x09))) | (x05 & x08 & ~x09 & ((x02 & ~x07) | (~x01 & ~x02 & x07)))) : ((x07 & x08 & x09 & x01 & x02 & x05) | (~x01 & ((x07 & ((x02 & ~x08 & (x05 ^ ~x09)) | (~x02 & ~x05 & x08 & x09))) | (~x02 & x05 & ~x07 & x08 & x09))))) : ((~x02 & ((x07 & ((~x01 & ((x00 & ~x08 & (x05 ^ ~x09)) | (x08 & ((~x05 & x09) | (~x00 & x05 & ~x09))))) | (~x00 & x01 & x05 & x08 & x09))) | (x01 & ~x07 & ((~x00 & ((x08 & ~x09) | (x05 & ~x08 & x09))) | (x08 & x09 & x00 & ~x05))))) | (~x00 & x01 & x02 & ~x05 & ~x07 & x08 & x09))))) | (~x06 & x07 & x08 & ~x09 & x10 & ~x02 & ~x05 & x00 & ~x01))) | (~x00 & ((~x02 & x05 & ((x01 & ~x06 & x09 & ((~x08 & x10 & ~x03 & x07) | (x08 & ~x10 & x03 & ~x07))) | (~x01 & x03 & x06 & x07 & x08 & ~x09 & ~x10))) | (x01 & x02 & ~x03 & ~x05 & x06 & ~x07 & ~x08 & ~x09 & ~x10))) | (x06 & x07 & ~x08 & ~x09 & ~x10 & x00 & x01 & ~x02 & ~x03 & x05);
endmodule