module pla__x9dn ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    z0, z1, z2, z3, z4, z5, z6  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26;
  output z0, z1, z2, z3, z4, z5, z6;
  assign z0 = x00 & x01 & x02 & x03 & x04 & x05 & ((x06 & ((~x07 & x08 & x09) | (~x08 & ~x09))) | (x07 & x13 & (x08 | x09)) | (~x07 & x10 & ~x11 & ~x12));
  assign z1 = ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & ((x07 & x16 & (x08 | x09)) | (~x07 & ((x08 & x09 & x14) | (~x11 & ~x12 & x15))) | (~x08 & ~x09 & x14));
  assign z2 = (((x06 & ((~x07 & x08 & x09) | (~x08 & ~x09))) | (x07 & x13 & (x08 | x09)) | (~x07 & x10 & ~x11 & ~x12)) & (~x17 | (x19 & (~x18 | (x21 & (~x20 | (~x22 & x23))))))) | (((x07 & x16 & (x08 | x09)) | (~x07 & ((x08 & x09 & x14) | (~x11 & ~x12 & x15))) | (~x08 & ~x09 & x14)) & (x17 | (~x19 & (x18 | (~x21 & (x20 | (x22 & ~x23)))))));
  assign z3 = (((x06 & ((~x07 & x08 & x09) | (~x08 & ~x09))) | (x07 & x13 & (x08 | x09)) | (~x07 & x10 & ~x11 & ~x12)) & (~x05 | (x04 & (~x03 | (~x01 & x02))))) | (((x07 & x16 & (x08 | x09)) | (~x07 & ((x08 & x09 & x14) | (~x11 & ~x12 & x15))) | (~x08 & ~x09 & x14)) & (x05 | (~x04 & (x03 | (x01 & ~x02)))));
  assign z4 = (~x24 | ~x25) & ((((~x07 & x08 & x09) | (~x08 & ~x09)) & ((x00 & x01 & x02 & x03 & x04 & x05 & x06 & x17 & x18 & x19 & x20 & x21 & x22 & x23 & x26) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x14 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26))) | (~x07 & ~x11 & ~x12 & ((x17 & x18 & x19 & x20 & x21 & x22 & x23 & x26 & x00 & x01 & x02 & x03 & x04 & x05 & x10) | (~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x15))) | (x07 & (x08 | x09) & ((x17 & x18 & x19 & x20 & x21 & x22 & x23 & x26 & x00 & x01 & x02 & x03 & x04 & x05 & x13) | (~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x16))));
  assign z5 = (((~x07 & x08 & x09) | (~x08 & ~x09)) & ((x00 & x01 & x02 & x03 & x04 & x05 & x06 & x17 & x18 & x19 & x20 & x21 & x22 & x23 & x26) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x14 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26))) | (~x07 & ~x11 & ~x12 & ((x17 & x18 & x19 & x20 & x21 & x22 & x23 & x26 & x00 & x01 & x02 & x03 & x04 & x05 & x10) | (~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x15))) | (x07 & (x08 | x09) & ((x17 & x18 & x19 & x20 & x21 & x22 & x23 & x26 & x00 & x01 & x02 & x03 & x04 & x05 & x13) | (~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & ~x23 & ~x26 & ~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x16)));
  assign z6 = (((~x07 & x08 & x09) | (~x08 & ~x09)) & ((x00 & x01 & x02 & x03 & x04 & x05 & x06 & x17) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x14 & ~x17))) | (~x07 & ~x11 & ~x12 & ((x00 & x01 & x02 & x03 & x04 & x05 & x10 & x17) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x15 & ~x17))) | (x07 & (x08 | x09) & ((x00 & x01 & x02 & x03 & x04 & x05 & x13 & x17) | (~x00 & ~x01 & ~x02 & ~x03 & ~x04 & ~x05 & x16 & ~x17)));
endmodule