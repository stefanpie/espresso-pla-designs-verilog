module pla__misex3 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n,
    r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  output r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2;
  assign r2 = ((k | (~j & l)) & ((b & ((f & ((~c & ((d & ~h & i & ~m & n) | (a & ~d & e & ~g & h & m & ~n))) | (~h & i & ~m & n & ((~e & (d | ~g)) | (~d & e & g))))) | (~g & h & m & ~n & ((a & ((c & ~d & e) | (d & ~e))) | (e & (~a | (~d & ~f))))) | (c & ~h & i & ~m & n & ((e & ~f) | (~d & ~e & g))))) | (c & ~h & i & ~m & ~n & ((f & (~d | ~e)) | (d & e & ~f))))) | (h & ((b & (m ? (~n & ((g & (l ? ~i : j)) | (k & ~l)) & ((e & (~a | (~d & (~f | (a & (c | (~c & f))))))) | (a & d & ~e))) : (n & (k ? (~i | ~j | ~l) : j) & ((c & ((e & ~f) | (~d & ~e & g))) | (f & ((d & (~c | ~e)) | (~d & e & g) | (~e & ~g))))))) | (c & ~m & ~n & ((f & (~d | ~e)) | (d & e & ~f)) & (k ? (~i | ~j | ~l) : j)))) | (b & g & m & ~n & ((e & (~a | (~d & (~f | (a & (c | (~c & f))))))) | (a & d & ~e)) & ((j & ((~i & (~k | l)) | (~k & l))) | (k & ((i & (~j | ~l)) | (~j & ~l))) | (~h & i & l)));
  assign s2 = ((k | (~j & l)) & ((c & ((~n & ((a & ~b & ~g & h & m & (e ? d : f)) | (d & ~h & i & ~m & (~e ^ ~f)))) | (~h & i & ~m & n & ((f & (~b | (~e & (~g | (b & (d | (~d & g))))))) | (b & e & ~f))))) | (d & ~n & ((~g & h & m & ((b & (a ^ e)) | (a & ~c & (~e | f)))) | (~c & f & ~h & i & ~m))))) | (h & ((~n & ((m & ((g & (l ? ~i : j)) | (k & ~l)) & ((d & ((b & (a ^ e)) | (a & ((~c & (~e | f)) | (~b & c & e))))) | (a & ~b & c & ~e & f))) | (d & ~m & (k ? (~i | ~j | ~l) : j) & (c ? (~e ^ ~f) : f)))) | (c & ~m & n & (k ? (~i | ~j | ~l) : j) & ((f & (~b | (~e & (~g | (b & (d | (~d & g))))))) | (b & e & ~f))))) | (g & m & ~n & ((j & ((~i & (~k | l)) | (~k & l))) | (k & ((i & (~j | ~l)) | (~j & ~l))) | (~h & i & l)) & ((d & ((b & (a ^ e)) | (a & ((~c & (~e | f)) | (~b & c & e))))) | (a & ~b & c & ~e & f)));
  assign t2 = ((k | (~j & l)) & ((f & ((~n & ((~g & h & m & ((b & (a ? (~c & ~d) : (~d | e))) | (a & ((c & ~d & e) | (d & (~b | ~e)))))) | (e & ~h & i & ~m & (c ^ d)))) | (e & ~h & i & ~m & n & (b ? (~c & d) : c)))) | (~h & i & ~m & ((e & ((~f & ((b & n & (c | ~d)) | (c & ~n))) | (b & ~d & g & n))) | (b & ~c & d & ~f & g & n))))) | (f & ((~n & ((m & ((b & (a ? (~c & ~d) : (~d | e))) | (a & ((c & ~d & e) | (d & (~b | ~e))))) & ((g & ((j & ((~i & (~k | l)) | (~k & l))) | (k & ((i & (~j | ~l)) | (~j & ~l))) | (~h & i & l) | (h & (l ? ~i : j)))) | (h & k & ~l))) | (e & h & ~m & (k ? (~i | ~j | ~l) : j) & (c ^ d)))) | (e & h & ~m & n & (k ? (~i | ~j | ~l) : j) & (b ? (~c & d) : c)))) | (h & ~m & (k ? (~i | ~j | ~l) : j) & ((e & ((~f & ((b & n & (c | ~d)) | (c & ~n))) | (b & ~d & g & n))) | (b & ~c & d & ~f & g & n)));
  assign u2 = ((~e | f) & ((i & (((k | (~j & l)) & ((~c & d & ~n & ((a & ~g & h & m) | (g & ~h & ~m))) | (~b & c & g & ~h & ~m & n))) | (a & ~c & d & g & m & ~n & ((j & (l ? ~k : h)) | (k & (~j | ~l)) | (~h & l))))) | (g & h & ~m & (k ? (~i | ~j | ~l) : j) & ((~b & c & n) | (~c & d & ~n))))) | (i & (((k | (~j & l)) & ((~n & ((~g & h & m & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((e & ((~d & ~f) | (c & (~d | ~f)))) | (f & ((d & ~e) | (~b & c))))))) | (c & g & ~h & ~m & (e ? (~f | (~d & f)) : f)))) | (b & g & ~h & ~m & n & (e ? (~c | ~f) : (d ? f : c))))) | (g & m & ~n & ((j & (l ? ~k : h)) | (k & (~j | ~l)) | (~h & l)) & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((e & ((~d & ~f) | (c & (~d | ~f)))) | (f & ((d & ~e) | (~b & c))))))))) | (g & h & ~m & (k ? (~i | ~j | ~l) : j) & ((c & ((~d & ((b & ~e & n) | (e & f & ~n))) | (~n & (~e ^ ~f)))) | (b & n & ((e & (~c | ~f)) | (d & ~e & f)))));
  assign n2 = (g & ((h & ((~n & ((m & ((j & ~k) | (~i & ~j & l)) & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f))))) | (~c & d & ~e & ~m & ((k & (~i | ~j)) | (i & j & ~k))))) | (~m & n & ((k & (~i | ~j)) | (i & j & ~k)) & ((c & (b ? ~d : ~e)) | (b & ((~c & d) | (e & (~d | ~f)))))))) | (k & m & ~n & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f)))) & ((i & (~h | ~j)) | (~j & ~l) | (~i & j & l))))) | (h & ~m & ((k & (~i | ~j)) | (i & j & ~k)) & ((~d & ((b & e & ~f & n) | (c & f & ~n))) | (c & ((e & ((b & ~g & n) | (~f & ~n))) | (f & (~g | (~b & n) | (~e & ~n))))) | (f & ((~c & d & ~n) | (b & n & ((~e & ~g) | (d & (~e | ~g))))))));
  assign o2 = h ? ((i & (j ? (~k & ~m & ((((~b & c & n) | (~c & d & ~n)) & (f | (~e & g))) | (b & n & ((c & (g ? ~d : e)) | (e & ((~d & (~f | g)) | (~f & g))) | (f & ((~e & ~g) | (d & (~e | ~g)))) | (~c & d & g))) | (c & ((f & (~g | (~n & (~d | ~e)))) | (e & ~f & ~n))))) : (k & ((g & ((~n & ((m & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f))))) | (~c & d & ~e & ~m))) | (~m & n & ((c & (b ? ~d : ~e)) | (b & ((~c & d) | (e & (~d | ~f)))))))) | (~m & ((~d & ((b & e & ~f & n) | (c & f & ~n))) | (c & ((e & ((b & ~g & n) | (~f & ~n))) | (f & (~g | (~b & n) | (~e & ~n))))) | (f & ((~c & d & ~n) | (b & n & ((~e & ~g) | (d & (~e | ~g)))))))))))) | (m & ~n & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f)))) & ((g & ((j & ~k) | (~i & ~j & k & l))) | (k & (~g | (~j & ~l)))))) : (i & k & ~m & ((((~b & c & n) | (~c & d & ~n)) & (f | (~e & g))) | (b & n & ((c & (g ? ~d : e)) | (e & ((~d & (~f | g)) | (~f & g))) | (f & ((~e & ~g) | (d & (~e | ~g)))) | (~c & d & g))) | (c & ((f & (~g | (~n & (~d | ~e)))) | (e & ~f & ~n)))));
  assign p2 = (~n & ((m & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f)))) & ((j & ((h & (g ^ k)) | (g & ((~i & (~k | l)) | (~h & i & k))))) | (g & ~h & i & ~k & l))) | (j & ~m & (h ? (~k | (~i & k)) : (i & k)) & (c ? (f ? (~d | ~e) : e) : (d & (f | (~e & g))))))) | (j & ~m & (h ? (~k | (~i & k)) : (i & k)) & ((n & ((c & (b ? (g ? ~d : e) : (f | (~e & g)))) | (b & ((e & ((~d & (~f | g)) | (~f & g))) | (f & ((~e & ~g) | (d & (~e | ~g)))) | (~c & d & g))))) | (c & f & ~g)));
  assign q2 = l & ((~n & (((~j | k) & ((~g & h & m & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f))))) | (~h & i & ~m & (c ? (f ? (~d | ~e) : e) : (d & (f | (~e & g))))))) | (g & (j ? ((m & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f)))) & (~h | ~k)) | (~c & d & ~e & h & ~m & (~k | (~i & k)))) : ((m & ((b & ((a & (f ? ~c : d)) | (e & ~f) | (~a & (e | (~d & f))))) | (a & ((d & ((~e & f) | (~c & (~e | f)))) | (e & ((~d & ~f) | (c & (~d | ~f)))) | (~b & c & f)))) & (i ? k : h)) | (~c & d & ~e & h & k & ~m)))) | (h & ~m & (j ? (~k | (~i & k)) : k) & (c ? (f ? (~d | ~e) : e) : (d & f))))) | (~m & ((n & ((c & (b ? (g ? ~d : e) : (f | (~e & g)))) | (b & ((e & ((~d & (~f | g)) | (~f & g))) | (f & ((~e & ~g) | (d & (~e | ~g)))) | (~c & d & g))))) | (c & f & ~g)) & (h ? (j ? (~k | (~i & k)) : k) : (i & (~j | k)))));
  assign h2 = ~n & ((g & ((l & ((e & ((~d & ((~c & f & ~m & ((~h & ~i & j & k) | (h & i & ~j & ~k))) | (a & c & m & ((~i & (h | j)) | (j & ~k) | (~h & i))))) | (c & m & ((~i & (h | j)) | (j & ~k) | (~h & i)) & (a ? ~f : b)))) | (c & m & ((~i & (h | j)) | (j & ~k) | (~h & i)) & ((b & (a ? (d & ~f) : (~d & f))) | (a & f & (~b | (d & ~e))))))) | (c & m & ((k & ((i & (~j | ~l)) | (~j & ~l))) | (j & ((h & ~l) | (~i & ~k)))) & ((b & (a ? (d & ~f) : (e | (~d & f)))) | (a & ((e & (~d | ~f)) | (f & (~b | (d & ~e))))))))) | (~g & ((h & ((c & m & (k | (~j & l)) & ((b & (a ? (d & ~f) : (e | (~d & f)))) | (a & ((e & (~d | ~f)) | (f & (~b | (d & ~e))))))) | (~c & ~d & ~f & i & j & k & l & ~m))) | (~c & ~d & ~f & ~h & ~i & ~k & ~l & ~m))) | (c & h & k & ~l & m & ((b & (a ? (d & ~f) : (e | (~d & f)))) | (a & ((e & (~d | ~f)) | (f & (~b | (d & ~e))))))));
  assign i2 = ((k | (~j & l)) & ((e & ((d & ((b & ~h & i & ~m & n & (g ? ~f : c)) | (~g & h & m & ~n & a & ~c & f))) | (a & ~g & h & m & ~n & ((~d & ~f) | (c & (~b | ~d)))))) | (b & ((~g & ((a & h & m & ~n & ((d & ~e) | (~c & ~d & f))) | (i & ~m & n & d & f & ~h))) | (d & ~h & i & ~m & n & ((~e & f) | (~c & g))))) | (~b & c & d & ~h & i & ~m & n & (f | (~e & g))))) | (~n & ((~d & ((~c & ((~m & ((~e & ~f & ~g & ((h & i & j & k & l) | (~h & ~i & ~k & ~l))) | (e & f & g & h & ~k & l & i & ~j))) | (a & b & f & m & ((g & ((j & ((~i & (~k | l)) | (~k & l))) | (k & ((i & (~j | ~l)) | (~j & ~l))) | (~h & i & l) | (h & (l ? ~i : j)))) | (h & k & ~l))))) | (a & e & m & (c | ~f) & ((g & ((j & ((~i & (~k | l)) | (~k & l))) | (k & ((i & (~j | ~l)) | (~j & ~l))) | (~h & i & l) | (h & (l ? ~i : j)))) | (h & k & ~l))))) | (g & ((d & (e ? ((~c & ((a & f & m & ((j & ((~i & (~k | l)) | (~k & l))) | (k & ((i & (~j | ~l)) | (~j & ~l))) | (~h & i & l) | (h & (l ? ~i : j)))) | (j & k & l & ~m & ~f & ~h & ~i))) | (c & f & ~h & ~i & j & ~k & ~l & ~m)) : ((l & ((c & ~f & ~m & ((~h & ~i & j & k) | (h & i & ~j & ~k))) | (a & b & m & ((~i & (h | j)) | (j & ~k) | (~h & i))))) | (a & b & m & ((k & ((i & (~j | ~l)) | (~j & ~l))) | (j & ((h & ~l) | (~i & ~k)))))))) | (a & ~b & c & e & m & ((j & ((~i & (~k | l)) | (~k & l))) | (k & ((i & (~j | ~l)) | (~j & ~l))) | (~h & i & l) | (h & (l ? ~i : j)))))) | (a & h & k & ~l & m & ((~b & c & e) | (d & ((b & ~e) | (~c & e & f))))))) | (d & ~m & n & (b ? ((g & ((~f & ((c & ~e & l & ((~h & ~i & j & k) | (h & i & ~j & ~k))) | (e & h & (k ? (~i | ~j | ~l) : j)))) | (~i & ((~c & h & k) | (c & e & f & ~k & ~l & ~h & j))) | (~c & h & (k ? (~j | ~l) : j)))) | (h & (k ? (~i | ~j | ~l) : j) & ((f & (~e | ~g)) | (c & e & ~g)))) : (c & ((h & (k ? (~i | ~j | ~l) : j) & (f | (~e & g))) | (e & ~f & g & ~h & k & l & ~i & j)))));
  assign j2 = (l & ((d & (c ? ((~e & ((b & ((h & i & ~k & ((~a & f & m & ~n & (g ^ j)) | (~f & g & ~j & ~m & n))) | (~f & g & ~h & ~i & ~m & n & j & k))) | (~f & g & ~m & ~n & ((~h & ~i & j & k) | (h & i & ~j & ~k))))) | (~b & e & ~f & g & i & ~k & ~m & n & (h ^ j))) : (e & ~f & g & i & ~k & ~m & ~n & (h ^ j)))) | (~c & ~d & j & k & ~m & ~n & ((~e & ~f & ~g & h & i) | (e & f & g & ~h & ~i))))) | (~c & ~d & ~f & ~g & ~h & ~i & ~j & ~k & ~l & ~m & ~n);
  assign k2 = (l & ((g & ((d & ((~m & (c ? ((h & i & ((((j & k & e & f) | (~j & ~k & ~e & ~f)) & (~n | (b & n))) | (~b & e & ~f & ~j & ~k & n))) | (~f & ~h & ~b & e & ~i & j & k & n)) : (e & ~f & ~n & ((~h & ~i & j & k) | (h & i & ~j & ~k))))) | (b & c & f & h & i & m & ~n & ((j & k & a & e) | (~j & ~k & ~a & ~e))))) | (~c & ~d & e & f & ~h & ~i & j & k & ~m & ~n))) | (~c & ~d & e & ~f & ~g & k & ~m & ~n & h & i & j))) | (~c & ~d & ~e & ~f & ~g & ~l & ~m & ~n & ~h & ~i & ~k);
  assign m2 = (l & (d ? (c ? ((h & ((i & ((b & ((f & ((m & ~n & ((~a & ~e & ~k & (g ^ j)) | (a & e & g & j & k))) | (e & g & j & k & ~m & n))) | (~e & ~f & g & ~m & n & ~j & ~k))) | (g & ~m & ((e & ((~j & ~k & n & ~b & ~f) | (f & j & k & ~n))) | (~e & ~f & ~j & ~k & ~n))))) | (~e & ~f & ~g & ~i & ~j & ~k & ~m & (~n | (~b & n))))) | (~f & g & ~h & j & ~m & ((n & ((~b & e & (i ^ k)) | (~i & k & b & ~e))) | (k & ~n & ~e & ~i)))) : (e & ~f & g & ~m & ~n & ((h & i & ~j & ~k) | (~h & j & (i ^ k))))) : (~n & ((~c & ~m & ((e & f & g & ((~h & ~i & j & k) | (h & i & ~j & ~k))) | (~f & ~g & h & i & j & k))) | (~a & b & c & ~e & ~f & g & ~h & ~i & ~j & k & m))))) | (~h & ~i & ~k & ~l & ~m & ((c & d & e & f & g & j & (~n | (b & n))) | (~c & ~d & ~f & ~g & ~n)));
  assign l2 = (~n & ((m & ((((a & b & c & (d ? (e & f) : ~e)) | (~e & ~f & (~a | ~d))) & (~k | ~l | (~g & (~j | k)))) | (d & ((~c & ((~b & e & ~f) | (~a & ~e))) | (~f & ((~a & ~e) | (~j & l & ~h & ~i))) | (~a & ~e & ((~g & (~j | k)) | ((~h | ~i) & (f | ~k)) | (f & k) | ~l | (g & j & ~k))) | (a & b & c & e & f & (~h | ~i | (~j & k))))) | (~e & ((~d & ((a & (~f | (b & c & f))) | (~f & (~b | ~c | h | i | j)))) | (h & ((~a & ~f) | (j & k & l & f & g & i))) | (~f & ((~b & c) | (~a & (~c | i | j)))))) | (~a & (~b | (f & g & h & i & j & k & l))) | ((a | e) & ((~j & ((g & h & i & ~k) | (~i & l & ~f & ~h))) | (~g & j & ~k))) | (~k & ((((~g & j) | (g & h & i & ~j)) & (~d | ~f | ~b | ~c)) | (~g & (~l | (~i & j))) | (~j & (~l | (~h & ~i & l))))) | (f & ((~j & l & ~h & ~i) | (~d & ((~b & ~c) | (j & k & l & g & h & i))))) | (l & (~b | ~c) & ((~h & ~i & ~j) | (g & h & i & j & k))) | (~h & (~g | (k & ~l & ~i & j))))) | (~m & ((d & ((k & ((c & e & f & g & ~i) | (~g & h & i & j & l))) | (~k & ((f & i & ((h & ~j) | (c & e & g & j))) | (~c & ~g & (h ? ~j : (j | ~l))))) | (~i & ((f & (c ? (e & g & (h | l)) : ~h)) | (~c & ~g & ~h))) | (c & e & f & g & (~j | (i & (~h | ~l)))))) | (~d & ((l & ((g & h & i & j & k) | (~c & ~g & ~i))) | (~c & ((h & (~i | (~f & g & j))) | ((f | g) & (i ? j : ~e)) | (~j & ((~e & (f | i)) | (g & ~i) | (i & (~f | ~g | ~h | k)))) | (f & (~g | (~h & i))) | (g & ((~f & (~i | (i & k))) | ~l | (~i & ~k))) | (~g & (i ? (~h | ~k) : k)) | (i & ~l))) | (c & ((~e & ~f & (~i | (i & ~j))) | (~i & (~h | (h & ~j & ~k))))) | (~f & ((h & i & ~j & ~k) | (g & ~h & ~i))) | (i & j & ~k & g & ~h))) | (~f & ((l & ((~c & ~g & ~i) | (i & j & k & c & h))) | ((c ^ e) & ((g & ((~i & (~j | ~k)) | (h & j) | (i & k))) | (i & ~j & (~h | k)))) | (~g & ((~h & (c ? ~e : i)) | (~i & (c ? (~e & k) : (h | k))) | (c & ~e & (i | j)) | (~c & i & (~j | ~k | ~l)))) | (c & ((~i & ((e & (~h | (h & ~j & ~k))) | (~h & ~l) | (~e & g & h))) | ((~l | (i & j)) & (~e | (~h & ~k))) | (~k & ~l & h & ~j))) | (g & ((~h & ~i & ~k) | (~c & e & ~l))) | (~c & e & (i ? ~l : h)))) | (~k & ((~j & ((h & ((c & ((e & (~g | i)) | (f & (i | (~i & l))) | (~g & ~l))) | (~e & (f | (~c & i))) | (f & ~g) | (~c & (~i | (g & ~l))))) | (~e & f & ~h & ~l))) | (~h & (g ? ((~c & (~i | ~l)) | (~e & i & j)) : ((i & j) | ((j | ~l) & (c | f))))))) | (g & ((~h & ~i & (~j | (~c & (~e | ~l)))) | (j & k & l & ~e & h & i))) | (l & ((c & ((f & ~h & ~i) | (~g & h & i & j & k))) | (~c & ((~g & ~h & ~i) | (i & j & k & f & h))) | (i & j & k & f & ~g & h))) | (~h & ~i & ((c & (~g | (f & k))) | (~g & (f | k)))))) | (i & ((j & k & l & ~f & g & h) | (~h & ~k & ~l))))) | (~m & ((n & ((~i & ((f & (((k | l) & (~h | (b & c & d & e & g))) | (b & c & d & e & g & h) | (~b & ~h))) | (~h & ((~f & (~l | (e & (b | ~k)))) | (~e & (~l | (g & (~b | ~k)))) | ~g | ~j | ~c | ~d)) | (~f & ((~b & e) | (b & c & d & ~e & g)) & (h | ~j | ~k)) | (~j & ~k & e & h))) | ((~c | ~d | ~e | ~f | ~g | (~b & f)) & ((h & i & j & k & l) | (~h & ~k & ~l))) | (~d & ((~f & ((~e & ~g) | (~b & (e | ~g)))) | (~c & (e ? (f & ~g) : g)) | (~k & (h ^ j)))) | (~k & (((h ^ j) & (~c | (~b & ~e & g))) | (~b & ((f & ~h & j) | (i & ~j & ~e & h))) | (~h & ((j & ((b & ~f & (e | i)) | ~g | (~e & (f | i)))) | (~l & (i | ~j)))) | (f & ((h & ~j) | (b & c & d & e & g & i))) | (h & ~j & ((b & (e | ~g)) | (e & ~g) | (~l & (~e | ~f)))))) | (~c & (~b | (~e & ~f & ~g))) | (~f & ((((~b & e) | (d & ~e & b & c)) & ((~j & (~h | k)) | (i & k) | ~l | (h & j))) | (~e & ((b & (~g | (i & j & c & d))) | (~g & (~h | i | j | k | ~l)))) | (~b & ~g & (j | k | ~l | e | ~h | i)))) | (b & c & d & e & f & g & (~j | (i & (~h | ~l)))))) | (f & ~h & (i ? (j & ~k) : ~e)) | (~g & ((h & i & ~j & ~k) | (~c & d & ~f))) | (h & ~j & ~k & (i ? ~l : g))));
endmodule