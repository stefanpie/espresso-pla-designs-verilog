module pla__in0 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10;
  assign z00 = (~x11 & ~x12 & ((~x01 & ((~x13 & ((~x10 & ((~x09 & (x00 ? (x03 | (x02 & ~x03)) : (x05 & (~x06 | (x06 & (x02 ? x07 : (~x07 | (x07 & (~x04 | (x03 & x04)))))))))) | (~x00 & x09 & (x02 | (~x02 & (x03 | (~x03 & (x04 | (~x04 & x05 & (~x06 | (x06 & ~x07))))))))))) | (x00 & ~x02 & ~x03 & x10 & x14))) | (x10 & (x00 ? x13 : (x14 | (x13 & ~x14)))))) | (x01 & (x10 ? (x14 | (x13 & ~x14)) : (~x13 & (x09 ? ~x00 : ((x02 & ((~x00 & ((~x05 & ((~x03 & (x04 ? ~x06 : (x06 & ~x07))) | (~x04 & (x06 ? x03 : ~x07)))) | (x03 & (x04 | (~x04 & ((x05 & (~x07 | (x06 & x07))) | (~x06 & x07))))))) | (x00 & (x03 ? (x05 ? ~x06 : x04) : (x05 ? ~x04 : ~x06))) | (~x03 & x04 & x05))) | (x00 & ((~x03 & ((~x02 & x04 & (x05 ? (x06 | (~x06 & ~x07)) : ~x06)) | (~x05 & x06))) | (~x04 & x05 & ~x02 & x03))) | (~x00 & ~x02)))))) | (x09 & ~x13 & (x10 ? ~x14 : x00)) | (~x09 & ~x10 & x13))) | (x09 & x10 & x11 & x12 & ~x13);
  assign z01 = ~x09 & ~x10 & ~x11 & ~x12 & ~x13 & (x01 ? ((x00 & ((x05 & (x02 ? (x03 ? x06 : ~x04) : (~x04 & x06))) | (~x02 & ~x04 & ~x05 & (x03 | (~x03 & ~x06))))) | (x02 & ~x03 & x04 & x05)) : (x00 ? (~x03 | (x02 & x03)) : (~x05 | (x05 & ~x06))));
  assign z02 = (x09 & x10 & x11 & x12 & ~x13) | (~x11 & ~x12 & ((~x09 & ~x10 & ((x03 & ((x00 & ~x01 & ~x13 & (~x04 | (x02 & x04))) | (~x02 & x13))) | (~x02 & ((~x03 & ~x04 & x13) | (~x00 & x01 & ~x13))) | (x02 & x13))) | (x10 & ((~x01 & (x00 ? (x13 | (~x02 & ~x03 & ~x13 & x14)) : (x14 | (x13 & ~x14)))) | (x01 & (x14 | (x13 & ~x14))) | (x09 & ~x13 & ~x14)))));
  assign z03 = ~x11 & ~x12 & (x13 ? x10 : ((~x00 & ~x01 & ~x02 & x05 & x06 & ~x09 & ~x10 & (~x07 | (x07 & (~x04 | (x03 & x04))))) | (x09 & x10 & ~x14)));
  assign z04 = (x09 & x10 & x11 & x12 & ~x13) | (~x11 & ~x12 & ((~x09 & ~x10 & ((~x13 & (x00 ? ((x02 & ((x01 & x03 & (x05 ? ~x06 : x04)) | (~x01 & ~x03 & x04 & ~x05 & ~x06))) | (~x01 & ~x02 & ~x03 & x05)) : (x01 ? ~x02 : (x05 & ~x06)))) | (~x02 & x13 & (x03 | (~x03 & ~x04))))) | (x10 & (x01 ? (x14 | (x13 & ~x14)) : (x00 ? (x13 | (~x02 & ~x03 & ~x13 & x14)) : (x14 | (x13 & ~x14)))))));
  assign z05 = ~x13 & ((~x10 & ~x11 & ~x12 & ((~x02 & ((x00 & x04 & ~x09 & ((x01 & ~x03 & x05 & (x06 | (~x06 & ~x07))) | (~x01 & x03 & ~x05 & x06 & ~x07))) | (~x00 & ~x01 & ~x03 & ~x04 & x05 & ~x06 & x09))) | (x01 & ~x09 & ((~x05 & ((x00 & ~x03 & (x06 | (x02 & ~x06))) | (~x00 & x02 & x03 & ~x04 & x06))) | (~x00 & x02 & x03 & (x04 | (~x04 & (x07 ? ~x06 : x05)))))))) | (~x09 & x10 & x11 & x12 & x14 & (~x02 ^ ~x03)));
  assign z06 = x12 ? (x10 ? (~x11 & x13) : x11) : (((x14 | (x13 & ~x14)) & (x11 | (x10 & ~x11 & (x00 ? x01 : (~x01 & ~x08))))) | (~x10 & ~x11 & (x09 ? (~x13 & (x00 | (~x00 & (x01 | (~x01 & (x02 | (~x02 & (x03 | (~x03 & (x04 | (~x04 & (~x05 | (x05 & x06 & x07))))))))))))) : ((~x03 & ((~x13 & ((x01 & ((x02 & (x00 ? (~x04 & x05) : (~x05 & (~x04 | (x04 & x06))))) | (x00 & ~x02 & ((~x05 & x06 & ~x07) | (~x04 & (~x06 | (x05 & x06))))))) | (x00 & ~x01 & (~x02 | (~x05 & ~x06 & x02 & x04))))) | (~x02 & ~x04 & x13 & (x00 ? x01 : (~x01 & ~x08))))) | (~x13 & (((~x05 | (x05 & ~x06)) & ((~x00 & ~x01) | (x00 & x01 & ~x02 & x03 & ~x04))) | (x00 & x03 & (x01 ? (x04 & (~x02 | (x02 & x05 & x06))) : x02))))))));
  assign z07 = (x01 & ((~x11 & ~x12 & ((~x09 & ~x10 & (x02 ? (x13 ? ~x00 : ((~x05 & (x00 ? (~x03 & (~x04 | (x04 & x06 & x07))) : (x03 & ~x04 & (x06 | (~x06 & ~x07))))) | (x03 & ((x04 & (~x00 | (x00 & x05 & x06))) | (~x00 & ~x04 & ((x05 & (~x07 | (x06 & x07))) | (~x06 & x07))))))) : ((~x00 & x13 & (x03 | (~x03 & ~x04))) | (x00 & x03 & ~x04 & ~x05 & ~x13)))) | (~x00 & x10 & (x14 | (~x14 & (x13 | (x09 & ~x13))))))) | (x11 & x12 & ~x13 & ~x00 & x09 & x10))) | (x12 & (~x10 | (x10 & ((~x11 & x13) | (~x00 & ~x01 & x08 & x09 & x11 & ~x13)))));
  assign z08 = (~x12 & (x11 ? (x14 | (x13 & ~x14)) : ((~x09 & ~x10 & (x13 ? (((x02 | (~x02 & x03)) & (x00 ? ~x01 : (x01 | (~x01 & x08)))) | (~x02 & ~x03 & ~x04)) : (x01 ? ((x02 & ((x03 & ((x04 & (~x00 | (x00 & x05 & x06))) | (~x00 & ~x04 & ((x05 & (~x07 | (x06 & x07))) | (~x06 & x07) | (~x05 & x06))))) | (~x03 & ((x00 & (~x05 | (~x04 & x05))) | (~x05 & x06 & ~x07 & ~x00 & ~x04))) | (~x00 & ~x04 & ~x05 & ~x06 & ~x07))) | (x00 & ~x02 & (x03 ? (~x04 & (~x05 | (x05 & ~x06))) : (~x05 & ~x07 & (x06 | (x04 & ~x06)))))) : (x00 ? ((x03 & (x02 | (~x05 & x06 & ~x07 & ~x02 & x04))) | (x02 & ~x03 & ~x05 & (~x04 | (x04 & ~x06)))) : (x05 & ~x06))))) | (x10 & (x01 ? (x14 | (~x14 & (x13 | (~x00 & x09 & ~x13)))) : ((~x00 & (x14 | (x13 & ~x14))) | (x00 & x13) | (~x13 & ((x00 & ((~x02 & ~x03 & x14) | (x09 & ~x14))) | (x09 & ~x14 & ~x00 & x08))))))))) | (x10 & x12 & ((~x11 & x13) | (x09 & x11 & ~x13 & (x00 ? ~x01 : (x01 | (~x01 & x08))))));
  assign z09 = (~x10 & ((~x09 & ~x11 & ~x12 & ((~x13 & (x00 ? ((x06 & ((x01 & (x02 ? ((x03 & ~x04 & x05) | (~x03 & x04 & ~x05 & ~x07)) : (~x03 & ((~x05 & ~x07) | (~x04 & x05 & x07))))) | (~x01 & ~x02 & x03 & x04 & ~x05 & ~x07))) | (~x01 & ((x02 & x04 & (x03 | (~x06 & x07 & ~x03 & ~x05))) | (~x02 & ~x03 & ~x04 & ~x05 & x07)))) : ((x01 & x02 & ~x03 & ~x04 & ~x05) | (~x06 & x07 & ~x01 & x05)))) | (~x02 & ~x03 & ~x04 & x13 & x14))) | (x12 & x13))) | (x13 & (x11 ? ~x12 : x10));
  assign z10 = (x14 & ((x10 & ~x11 & (x12 ? x13 : (~x13 & (x01 | (~x01 & (~x00 | (x00 & ~x02 & ~x03))))))) | (x11 & ~x12) | (~x10 & x12))) | (~x11 & ~x12 & ((x13 & ~x14 & (x10 | (~x02 & ~x03 & ~x04 & ~x09 & ~x10))) | (~x09 & ~x10 & ~x13 & ((~x04 & ((x01 & ((~x03 & ((x02 & (x00 ? x05 : (~x05 & (~x06 ^ ~x07)))) | (x00 & ~x02 & (x05 ^ ~x06)))) | (x00 & x03 & x05 & (x02 ? (x06 & x07) : ~x06)))) | (x00 & ~x01 & (x02 ? x03 : (~x03 & ~x05 & (~x07 | (~x06 & x07))))))) | (x00 & x04 & ((x01 & ((x02 & x03 & x05 & x06) | (~x02 & ~x03 & ~x05 & ~x07))) | (~x05 & ~x06 & ~x07 & ~x01 & x02 & ~x03))) | (~x00 & ~x01 & x05 & ~x06 & ~x07)))));
endmodule