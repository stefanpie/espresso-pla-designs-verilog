module pla__cps ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23,
    z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010, z011,
    z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022, z023,
    z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034, z035,
    z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046, z047,
    z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058, z059,
    z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070, z071,
    z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082, z083,
    z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094, z095,
    z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106, z107,
    z108  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23;
  output z000, z001, z002, z003, z004, z005, z006, z007, z008, z009, z010,
    z011, z012, z013, z014, z015, z016, z017, z018, z019, z020, z021, z022,
    z023, z024, z025, z026, z027, z028, z029, z030, z031, z032, z033, z034,
    z035, z036, z037, z038, z039, z040, z041, z042, z043, z044, z045, z046,
    z047, z048, z049, z050, z051, z052, z053, z054, z055, z056, z057, z058,
    z059, z060, z061, z062, z063, z064, z065, z066, z067, z068, z069, z070,
    z071, z072, z073, z074, z075, z076, z077, z078, z079, z080, z081, z082,
    z083, z084, z085, z086, z087, z088, z089, z090, z091, z092, z093, z094,
    z095, z096, z097, z098, z099, z100, z101, z102, z103, z104, z105, z106,
    z107, z108;
  assign z000 = ~x04 & ((x09 & (x07 ? ((x08 & ((x10 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ((x01 & ((~x22 & ((x17 & x19 & (x20 | x21)) | (~x20 & ~x21 & ~x17 & ~x19))) | (~x17 & ~x19 & x20 & x21 & x22 & (x00 ? (x02 & x03) : (~x02 & ~x03))))) | (~x01 & x17 & x19 & x20 & x22))) | ~x11 | ~x12)) | (~x06 & ~x08 & x10 & x12)) : (x11 & (x08 ? (~x10 & x12) : x10)))) | (x07 & ~x08 & ((x11 & ((x10 & x12) | (~x09 & (x10 | x12)))) | (~x09 & ~x11 & ~x12))));
  assign z001 = ~x04 & ((~x08 & ((x11 & ((~x07 & x09 & (x10 | (~x10 & x12))) | (~x09 & ~x10 & x12) | (x10 & ~x12))) | (x07 & (~x09 | ~x10 | ~x11)))) | (x07 & ((~x09 & (x10 | x11)) | (~x11 & (x09 | x10)) | ~x12 | (x08 & x10 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x20 & (x18 ? ((~x17 & x19 & (x01 ? (~x21 | x22) : x21)) | (~x01 & x17 & ~x19 & x21 & ~x22)) : ((~x22 & ((x01 & (x17 ? (x19 & x21) : ~x19)) | (~x17 & ~x19 & x21))) | (x01 & ~x17 & ~x19 & ~x21)))) | (~x17 & ((x20 & (x18 ? ((~x01 & (~x19 | ~x21)) | (~x21 & (~x19 | ~x22))) : (~x19 & x21 & (x01 | x22)))) | (~x01 & x18 & ~x21 & ~x22))))))));
  assign z002 = ~x04 & ((x07 & ((x11 & (x08 ? (x10 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x17 & ((x21 & ((~x19 & x20 & ((~x01 & (x18 | (x02 & x22))) | (~x18 & ((x01 & (x03 ? (~x00 | ~x02) : x00)) | (x02 & ~x03 & x22))))) | (~x18 & ~x22 & (x01 | ~x20)) | (~x01 & x18 & x19 & ~x20))) | (~x20 & (x01 ? ((x18 & x19 & (~x21 | x22)) | (~x18 & ~x19 & ~x21 & x22)) : (~x22 & (x19 | (x18 & ~x21))))) | (~x18 & x19 & ~x22))) | (~x01 & ~x22 & ((~x18 & x19 & x20) | (x17 & x18 & ~x19 & ~x20 & x21))))) : (~x10 & ~x12))) | (~x08 & x09 & (~x10 | ~x12 | (x06 & ~x11))))) | (~x07 & ((x08 & (~x11 | ~x12)) | (~x10 & (x09 ? (~x11 | (~x08 & x11 & x12)) : x11)) | (~x09 & (x12 | (x10 & ~x11))))) | (~x09 & (x08 | (~x11 & x12))));
  assign z003 = ~x12 & ~x11 & x10 & x09 & x08 & ~x04 & x07;
  assign z004 = ~x12 & ~x11 & ~x10 & x09 & x08 & ~x04 & x07;
  assign z005 = x12 & ~x11 & x10 & x09 & ~x08 & ~x04 & x07;
  assign z006 = ~x12 & x11 & x10 & ~x09 & ~x08 & ~x04 & ~x07;
  assign z007 = ~x22 & x21 & ~x20 & ~x19 & x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z008 = x22 & ~x21 & ~x20 & ~x19 & x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z009 = x22 & ~x21 & ~x20 & ~x19 & x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z010 = ~x22 & ~x21 & ~x20 & ~x19 & x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z011 = ~x22 & ~x21 & ~x20 & ~x19 & x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z012 = ~x22 & x21 & ~x20 & x19 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z013 = x22 & x21 & x20 & x19 & x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z014 = ~x22 & x21 & ~x20 & x19 & x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z015 = ~x22 & ~x21 & ~x20 & x19 & x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z016 = x22 & x21 & x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z017 = ~x22 & x21 & x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z018 = ~x22 & x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z019 = ~x22 & x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z020 = x22 & ~x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z021 = ~x22 & ~x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z022 = ~x22 & ~x21 & ~x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z023 = (x08 & (~x10 | ~x11)) | (~x11 & (x09 ? (x10 & x12) : ~x12)) | x04 | ~x07 | (x11 & ((~x09 & (x10 | x12)) | (x10 & (x01 | ~x08 | ~x12 | x13 | x14 | x15 | x16 | x17 | ~x18 | ~x21 | x22 | x19 | ~x20))));
  assign z024 = ~x04 & ((~x07 & ((~x05 & ((x08 & (~x09 | ~x12)) | (~x10 & ((x09 & ~x11) | (~x08 & x12))) | (~x09 & (x10 | x11 | x12)))) | (x10 & x11 & ~x08 & x09))) | (x07 & ((x09 & ~x12 & (x08 | (x10 & x11))) | (x08 & ((~x09 & (x10 | x12)) | ~x11 | (x10 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x01 & (x17 ? ((~x18 & x19 & x20) | (~x05 & x18 & ~x19 & ~x20 & x21 & ~x22)) : ((~x05 & ((~x18 & x19) | (~x21 & ~x22 & x18 & ~x20))) | (x18 & ((x19 & (x20 ? (~x21 | x22) : (x21 | ~x22))) | (x20 & x21 & x22)))))) | (~x18 & ((~x22 & ((x19 & (x17 ? (x20 | (x01 & x21)) : ~x05)) | (x01 & ~x17 & ~x19 & (x20 ^ ~x21)))) | (~x05 & ~x17 & ((x19 & ~x20) | (~x21 & x22 & x01 & ~x19))))) | (~x17 & x18 & x19 & ((x01 & ~x20 & (~x21 | x22)) | (x20 & ~x21 & ~x22))))))))) | (~x05 & ((~x09 & x10 & x11) | (x08 & ~x11))));
  assign z025 = ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & x20 & x21 & x22 & ((x02 & ~x03 & (~x00 | ~x01)) | (x00 & x01 & ~x02 & x03));
  assign z026 = ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x18 & ~x19 & x20 & x21 & x22 & ((x03 & (~x00 | ~x01)) | (x00 & x01 & ~x03));
  assign z027 = ~x04 & x05 & ((x11 & (x09 ? (x12 & (x07 ? (x08 & x10 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x19 & ~x20 & ((~x01 & x18 & ~x22 & (~x17 ^ x21)) | (x01 & ~x17 & ~x18 & ~x21 & x22))) | (x19 & ~x22 & ~x17 & ~x18))) : (~x08 & ~x10))) : (~x07 | (~x08 & x10)))) | (~x07 & ((x08 & (~x11 | ~x12)) | (~x09 & (x10 | x12)) | (x09 & ~x10 & ~x11))));
  assign z028 = ~x04 & (((~x11 | ~x12) & (x07 ? (~x08 & x09) : x08)) | (~x08 & ~x10 & (x07 ? (x09 | (x11 & ~x12)) : x12)) | (~x09 & ((x08 & (x11 | ~x12)) | (x11 & ~x12 & ~x07 & x10))));
  assign z029 = ~x04 & ((x12 & ((x07 & ~x08 & (x09 ? (x10 & x11) : ~x10)) | (~x07 & x08 & x09 & ~x10 & x11))) | (x07 & ~x08 & ~x09 & ~x10 & ~x11));
  assign z030 = ~x04 & x07 & ((x08 & x09 & ~x10 & (x11 ^ x12)) | (x10 & x11 & ~x08 & ~x09));
  assign z031 = ~x04 & ((x10 & (x07 ? (x08 & x09 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ((~x01 & ((x18 & ((~x21 & ~x22) | (~x19 & x20))) | (x19 & (~x21 | x22 | ~x18 | ~x20)))) | (~x21 & (x19 ? (x20 & ~x22) : ((x18 & x20) | (x01 & ~x18 & x22)))) | (~x18 & ((~x20 & x21 & ~x22) | (x19 & (~x20 | ~x22)))) | (x19 & ~x20 & x22))) : (~x08 & ~x09 & (~x11 | x12)))) | (~x10 & ~x11 & ~x12 & ~x07 & ~x08 & x09));
  assign z032 = ~x22 & x20 & x19 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z033 = ~x04 & x07 & ((x08 & ((x10 & ((x12 & (~x09 | (x11 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x17 & ((x21 & ((x00 & ((x18 & x19 & ~x20) | (x01 & ~x18 & ~x19 & ~x22))) | (~x20 & ((x01 & (x18 ? x19 : (~x19 & ~x22))) | (x18 & x19 & ~x22))) | (~x01 & ~x19 & x20 & x22 & (x02 | x18)))) | (x19 & ~x20 & x22 & x01 & x18))) | (~x01 & x17 & ~x18 & ~x21 & ~x22 & x19 & x20))))) | (~x09 & (x00 | ~x11)))) | (~x09 & x11 & (x00 | x12)))) | (~x08 & x09 & x10 & x11 & ~x12));
  assign z034 = ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x21 & ((~x01 & x02 & ~x18 & ~x19 & x20 & x22) | (x01 & x18 & x19 & ~x20 & ~x22));
  assign z035 = ~x04 & x07 & x08 & ((x10 & (x09 ? (x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ((~x20 & ((x01 & ((~x21 & x22 & x18 & x19) | (x21 & ~x22 & ~x18 & ~x19))) | (x18 & x19 & x21 & (~x01 | ~x22)))) | (x02 & ~x18 & ~x19 & x20 & x21 & x22 & (~x00 | ~x01 | ~x03)))) : (~x11 | ~x12))) | (x11 & x12 & ~x09 & ~x10));
  assign z036 = ~x04 & x07 & x10 & x11 & (x08 ? (x12 & (~x09 | (~x13 & ~x14 & ~x15 & ~x16 & ((~x01 & x20 & ((~x17 & x18 & ~x19 & x21 & x22) | (x17 & ~x18 & x19 & ~x21 & ~x22))) | (x01 & ~x17 & x18 & x19 & ~x20 & x21 & x22))))) : (x09 & ~x12));
  assign z037 = ~x04 & ((x08 & ((x07 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x17 & ((~x22 & ((~x20 & ((~x01 & (~x18 ^ ~x21)) | (x19 & ~x21))) | (~x18 & (x19 | (x20 & x21 & ~x00 & x01))))) | (x01 & ~x18 & ~x19 & x22 & ((~x20 & ~x21) | (~x02 & x20 & x21 & (x00 | x03)))))) | (~x01 & x21 & ~x22 & ((~x18 & x19 & x20) | (x17 & x18 & ~x19 & ~x20))))) | ((~x11 | ~x12) & (~x07 | (~x09 & ~x10))))) | (x09 & ((~x07 & ~x10 & (~x11 | (~x08 & x11 & x12))) | (x06 & x07 & ~x08 & x10 & ~x11 & x12))) | (~x07 & ~x09 & (x10 | x11 | x12)));
  assign z038 = ~x04 & ((x07 & ((x09 & ((~x06 & ~x08 & x10 & x12) | (x08 & ~x11))) | (~x08 & ((x10 & x11) | (~x09 & (~x11 ^ x12)))) | (x10 & ((~x09 & (x08 | ~x12)) | (x08 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & (x17 ? (~x18 & x19 & (x01 ? (~x22 & (x20 | x21)) : (x20 & (~x21 | x22)))) : ((x21 & ((~x01 & ((x18 & x19 & ~x20) | (~x02 & x03 & ~x19 & x20 & x22))) | (x01 & ~x18 & ~x19 & ((x20 & x22 & (x02 | (~x00 & ~x03))) | (x00 & ~x22))) | (~x20 & x22 & x18 & x19))) | (x18 & x20 & ((~x21 & ~x22) | (~x19 & (~x21 | (~x01 & x22))))) | (x01 & ~x18 & ~x19 & ~x20 & ~x22)))))))) | (x09 & x11 & ((~x08 & x10) | (~x10 & x12 & ~x07 & x08))));
  assign z039 = ~x04 & ((x09 & ((x07 & ((x08 & x10 & x11 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x17 & ((~x18 & ((x21 & ((x20 & ((x01 & ((x00 & ~x02 & ~x19 & x22) | (~x00 & ~x22))) | (~x02 & x03 & ~x19 & x22))) | (~x01 & ~x20 & ~x22))) | (x19 & ~x22) | (x01 & ~x20 & ~x21 & (~x19 | ~x22)))) | (~x21 & (x01 ? (x19 & ~x22) : (x18 & ((x19 & x20 & x22) | (~x20 & ~x22))))) | (~x01 & x18 & ~x19 & x20 & x21 & ~x22))) | (~x18 & x19 & ((~x22 & ((x20 & x21) | (x01 & (x20 | x21)))) | (~x01 & x17 & x20 & x22))) | (~x01 & x17 & x18 & x21 & ~x22 & ~x19 & ~x20))) | (~x11 & x12) | (~x08 & (~x10 | ~x11)))) | (x08 & (x11 ? ~x12 : ~x07)) | (~x07 & ((~x10 & ~x11) | (~x08 & x11 & (x10 | (~x10 & x12))))))) | (x07 & ((~x08 & x12 & (~x11 | (~x09 & x10))) | (~x10 & x11 & ~x12))) | (~x09 & ((x08 & (x11 ? ~x07 : ~x10)) | (~x07 & (x11 ? (~x10 | ~x12) : x10)))) | (~x07 & x08 & x11 & ~x12));
  assign z040 = ~x04 & ((x08 & ((~x09 & (~x07 | (~x10 & ~x11))) | (~x10 & (~x07 | (x11 & ~x12))) | (~x07 & (~x11 | ~x12)) | (x09 & (x11 ? (~x12 | (x07 & x10 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x01 & x21 & ~x22 & ((~x18 & x19 & x20) | (x17 & x18 & ~x19 & ~x20))) | (~x17 & ((~x22 & ((x19 & (~x18 | (x01 & ~x20))) | (x20 & (x01 ? ((x18 & ~x21) | (~x00 & ~x18 & x21)) : (x18 & ~x19))) | (~x01 & ~x20 & (~x18 ^ ~x21)))) | (x20 & ((x22 & ((~x18 & ~x19 & x21 & (x01 ? (~x02 | (x00 & x03)) : x02)) | (~x01 & x18 & ~x21))) | (~x19 & ~x21 & x01 & x18))) | (x01 & ~x18 & ~x19 & ~x20 & ~x21 & x22)))))) : x12)))) | (~x08 & ((~x10 & ((x09 & (x07 | (~x07 & x11 & x12))) | (~x11 & x12) | (x07 & (~x11 | ~x12)))) | (x07 & ((~x11 & (x06 | ~x09 | ~x12)) | (x10 & x11 & x12))))) | (~x07 & ~x09 & (x11 | (x10 & x12))));
  assign z041 = ~x04 & x07 & ((~x08 & x09 & x10 & x11 & ~x12) | (x08 & ((x10 & (~x09 | (x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x01 & x17 & ~x18 & ~x21 & ~x22 & x19 & x20) | (~x17 & ((~x20 & ((x01 & ((x21 & ~x22 & ~x18 & ~x19) | (x18 & x19 & x22))) | (x18 & x19 & x21))) | (~x19 & x20 & x21 & x22 & ((~x01 & (x02 | x18)) | (x02 & ~x18 & (~x00 | ~x03)))))))))) | (~x09 & x11 & x12))));
  assign z042 = ~x04 & ((x10 & ((x08 & ~x11) | (x07 & ((~x08 & (x09 ? x12 : x11)) | (x09 & (~x11 | (x08 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x01 & (x17 ? ((~x18 & x19 & x20) | (x18 & ~x19 & ~x20 & x21 & ~x22)) : (x18 & ((x21 & ~x22 & ~x19 & x20) | (x19 & (x20 ^ x21)))))) | (~x17 & ((~x18 & ((~x19 & ((x20 & x21 & x22) | (x01 & (x20 ^ ~x21)))) | (~x22 & (x19 | (~x20 & (x01 | x21)))))) | (x19 & ((~x21 & ~x22) | (~x20 & (~x22 | (x01 & x18 & ~x21))))))) | (~x18 & x19 & x20 & ~x22))))))))) | (~x07 & ((~x09 & (x08 | x12)) | (x08 & (~x10 | ~x11)) | (~x10 & ~x11 & x12))) | (x08 & ((~x09 & ~x10 & x11) | ~x12 | (x09 & ~x11))));
  assign z043 = ~x04 & x07 & ((~x08 & ~x09 & ~x10 & (~x11 | ~x12)) | (~x01 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x17 & x18 & ~x15 & ~x16 & ~x21 & ~x22 & ~x19 & ~x20));
  assign z044 = ~x04 & ((x09 & ((~x08 & x11 & x12 & (~x07 ^ x10)) | (~x11 & (x08 | (x07 & x10 & ~x12))) | (x07 & x08 & x10 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x17 & ((~x18 & ((~x19 & (x20 ? (x21 & (x01 | x22)) : (~x21 & x22))) | (~x22 & (x19 | (~x20 & x21))))) | (~x01 & x18 & ((x21 & ~x22 & ~x19 & x20) | (~x20 & (x21 ? x19 : ~x22)))) | (x19 & ~x22 & (~x20 | ~x21)))) | (~x18 & x19 & x20 & ~x22) | (~x01 & x17 & (x18 ? (~x19 & ~x20 & (~x21 | ~x22)) : (x19 & x20))))))) | (~x09 & (x07 ? (~x10 & (~x12 | (~x08 & ~x11))) : (x08 | x12))) | (~x07 & ((x08 & (~x10 | ~x11)) | (~x10 & ~x11 & x12))) | (x08 & (~x12 | (x10 & ~x11))));
  assign z045 = ~x04 & x09 & x10 & (x07 ? (x08 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ((x17 & ((~x19 & ((x21 & x22) | (~x01 & (~x20 | x21)))) | (~x20 & (x22 | (x01 & x19 & x21))))) | (~x01 & ~x19 & ~x20 & ~x21 & ~x22))) : ~x08);
  assign z046 = ~x04 & x07 & x08 & x11 & x12 & ((~x09 & ~x10) | (~x13 & ~x14 & ~x15 & x01 & x09 & x10 & ~x16 & ~x17 & x18 & x19 & ~x20 & ~x21 & x22));
  assign z047 = ~x04 & x12 & ((x09 & x11 & ((x01 & (x07 ? (~x08 & x10) : (x08 & ~x10))) | (x07 & x08 & x10 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x18 & x19 & ~x20))) | (~x07 & ~x09 & ((~x10 & ~x11) | (x01 & ~x08 & x10))));
  assign z048 = x22 & x20 & x19 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z049 = ~x22 & x20 & x19 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z050 = ~x04 & (x07 ? (x09 & x10 & x11 & x12 & (~x08 | (~x13 & ~x14 & ~x15 & ~x16 & ~x18 & x19 & ((x20 & (~x22 | (~x01 & x17))) | (~x17 & ~x22))))) : ((~x09 & (x08 | (x10 & x12))) | (x08 & (~x10 | ~x11 | ~x12))));
  assign z051 = ~x04 & ~x07 & x08 & ((~x11 & ~x12) | (~x09 & x11 & x12));
  assign z052 = ~x04 & x12 & ((x10 & ((x01 & ~x08 & (x07 ? (x09 & x11) : ~x09)) | (x07 & x08 & x09 & x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x20 & ((~x17 & ~x18 & x19) | (~x19 & x21 & ~x22 & ~x01 & x17 & x18))))) | (~x07 & ~x10 & ((x09 & x11 & x01 & x08) | (~x09 & ~x11))));
  assign z053 = ~x04 & (x07 ? (x09 & x10 & x11 & x12 & (~x08 | (~x13 & ~x14 & ~x15 & ~x16 & ~x18 & x19 & ((x20 & (~x22 | (~x01 & x17))) | (~x17 & ~x22))))) : ((~x09 & (x08 | (x10 & x12))) | (x08 & (~x11 | ~x12)) | (~x10 & (x08 | (~x11 & x12)))));
  assign z054 = ~x04 & ((x08 & (x07 ? (x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ((~x18 & x19 & x20 & ~x22) | (~x01 & ((~x18 & x19 & x20) | (x18 & ~x19 & ~x20 & x21 & ~x22))))) : (~x09 | ~x11 | ~x12))) | (~x11 & x12 & ~x07 & ~x10));
  assign z055 = ~x04 & x09 & x10 & (x07 ? (x08 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ((x20 & ((x19 & ~x22) | (~x01 & (x19 | x21)))) | (x21 & ~x22 & x01 & x19))) : (~x08 & ~x12));
  assign z056 = ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & x21 & ((~x19 & (~x01 | x22)) | (~x01 & (x20 | x22)) | (~x20 & (x22 | (x01 & x19))));
  assign z057 = ~x04 & x09 & x10 & (x07 ? (x08 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ((x20 & ((x19 & ~x22) | (~x01 & (x19 | x21)))) | (x01 & ((~x20 & x22) | (x21 & (~x19 ^ ~x22)))))) : ~x08);
  assign z058 = x21 & x20 & ~x19 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z059 = ~x04 & ((x09 & (x07 ? (x08 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x17 & ~x18 & x19 & x20 & (~x01 | ~x22)) | (~x21 & ~x22 & ~x19 & ~x20 & x01 & x17 & x18))) : ((x08 & (~x11 | ~x12)) | (~x10 & (x08 | (~x11 & x12)))))) | (~x07 & ~x08 & ~x09 & x10 & x12));
  assign z060 = ~x01 & ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ~x20 & ~x21 & (~x19 | x22);
  assign z061 = ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & x19 & x20 & ~x21 & (~x01 | ~x22);
  assign z062 = x22 & ~x21 & ~x20 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z063 = ~x01 & ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ~x20 & x21 & (~x19 | x22);
  assign z064 = x01 & ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & x21 & x22 & (~x19 | ~x20);
  assign z065 = ~x04 & ((~x07 & ~x08 & ~x09 & x10 & x12) | (x09 & ((x12 & (x07 ? (x10 & x11 & (~x08 | (~x13 & ~x14 & ~x15 & ~x16 & ~x18 & x19 & x20 & ((~x01 & (~x17 | x22)) | (~x22 & (x01 | ~x17)))))) : (~x10 & ~x11))) | (~x07 & x08 & (~x10 | ~x11 | ~x12)))));
  assign z066 = ~x04 & ((x09 & ((x08 & (x07 ? (x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x21 & ~x22 & ~x19 & ~x20 & x01 & x17 & x18) | (~x18 & ((x20 & ((x19 & ~x22) | (~x01 & (x19 | (x17 & x21))))) | (x01 & x17 & ((~x20 & x22) | (x21 & (~x19 ^ ~x22)))))))) : (~x10 | ~x11 | ~x12))) | (~x07 & ((~x08 & x10) | (~x11 & x12))))) | (x10 & x12 & ~x07 & ~x08));
  assign z067 = ~x01 & ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ~x20 & (~x19 | x22);
  assign z068 = ~x04 & x09 & x10 & x11 & ((~x07 & ~x08) | (x01 & x07 & x08 & ~x14 & ~x15 & x12 & ~x13 & ~x16 & x17 & ~x18 & x21 & ~x22 & x19 & ~x20));
  assign z069 = ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ((x17 & x19 & (~x20 ^ ~x22)) | (~x20 & ~x21 & ~x22 & ~x01 & ~x17 & ~x19));
  assign z070 = ~x04 & x08 & x09 & (x07 ? (x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & ((~x01 & (x17 ? (~x19 & ~x20) : (x19 & x20))) | (~x20 & x22 & x17 & ~x19))) : ~x12);
  assign z071 = x21 & x20 & ~x19 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & ~x04 & x07;
  assign z072 = ~x04 & x10 & ((x08 & (x07 ? (x09 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x18 & x19 & ((~x01 & (x17 ? (x20 & ~x22) : x21)) | (~x17 & x21 & (~x20 | ~x22)))) : (~x11 | ~x12))) | (~x07 & ~x09 & (~x11 ^ x12)));
  assign z073 = ~x04 & ((x07 & ((~x09 & ~x10 & x11 & (x08 | ~x12)) | (x08 & (((~x11 | ~x12) & (x09 | x10)) | (x09 & x10 & ~x13 & ~x14 & ~x15 & ~x16 & ((~x17 & ((~x19 & ((~x18 & (x20 ? (x21 & (x01 | x22)) : ((~x01 & (~x21 | ~x22)) | (x21 & ~x22) | (~x21 & x22)))) | (~x01 & x18 & x20 & x21 & ~x22))) | (x18 & ((x19 & (x20 ? (~x21 & (~x01 | ~x22)) : (x01 ? (~x21 | ~x22) : x21))) | (~x21 & ~x22 & ~x01 & ~x20))))) | (~x01 & x17 & x18 & ~x19 & ~x20 & ~x21))))))) | (~x07 & ~x08 & ~x10 & x11 & x12));
  assign z074 = ~x04 & x07 & x10 & x11 & (x08 ? (x12 & (~x09 | (~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & x21 & x22 & (x01 ? (x19 & ~x20) : (~x19 & x20))))) : (x09 & ~x12));
  assign z075 = ~x04 & x09 & x10 & (x07 ? (x08 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & x17 & ~x18 & ((~x19 & ((x21 & x22) | (~x01 & (~x20 | x21)))) | (~x20 & (x22 | (x01 & x19 & x21))))) : ~x08);
  assign z076 = x22 & x21 & x20 & ~x19 & ~x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & ~x04 & x07;
  assign z077 = ~x04 & x07 & x08 & ((x09 & x10 & x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & x19 & ((~x22 & (~x20 | ~x21)) | (~x01 & (x20 ^ x21)))) | ~x12 | (~x09 & ~x11));
  assign z078 = ~x04 & x07 & x08 & (x09 ? (x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ((x21 & ((~x01 & ((x18 & x19 & (~x20 | x22)) | (~x18 & ~x19 & ~x20 & ~x22))) | (~x18 & ~x19 & x20 & (x01 | x22)))) | (x18 & x19 & ~x20 & ~x21 & ~x22))) : (~x11 | ~x12));
  assign z079 = ~x04 & x07 & x08 & (x09 ? (x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & x19 & ~x20 & (~x22 | (~x01 & x21))) : (~x11 | ~x12));
  assign z080 = ~x04 & x07 & x08 & (x09 ? (x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ((x18 & x19 & ~x20 & (~x22 | (~x01 & x21))) | (x20 & x21 & ~x22 & x01 & ~x18 & ~x19))) : (~x11 | ~x12));
  assign z081 = ~x04 & x07 & x08 & (x09 ? (x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & x19 & ~x20 & (~x22 | (~x01 & x21))) : (~x12 | (~x10 & ~x11)));
  assign z082 = ~x04 & x07 & x08 & ((~x09 & (x10 | ~x11)) | ~x12 | (x10 & x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & x19 & ((~x20 & (x21 | ~x22)) | (~x21 & (~x22 | (~x01 & x20))))));
  assign z083 = ~x04 & x07 & x08 & (x09 ? (x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & ~x20 & ((~x01 & x21 & (x18 ? x19 : (~x19 & ~x22))) | (~x21 & ~x22 & x18 & x19))) : (~x11 | ~x12));
  assign z084 = ~x04 & x07 & x08 & x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ((x22 & ((~x01 & ((x17 & ~x18 & ~x19) | (~x17 & x18 & x19 & x20 & x21))) | (x17 & ~x18 & (~x20 | (~x19 & x21))))) | (x19 & x20 & ~x22 & x17 & ~x18));
  assign z085 = ~x11 & ~x10 & ~x09 & ~x08 & ~x04 & x07;
  assign z086 = ~x04 & x07 & ((x09 & ((x12 & (x08 ? (x10 & x11 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & ~x19 & x20 & ~x22 & (x01 | ~x21)) : ~x11)) | (~x08 & ~x10 & ~x11))) | (~x08 & ~x09 & (x10 ? ~x11 : (x11 & x12))));
  assign z087 = ~x04 & x07 & (x08 ? (x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & ~x19 & ((~x21 & ~x22 & ~x01 & ~x20) | (x20 & x22 & (x01 | ~x21)))) : ((~x09 & ~x10 & (~x11 | ~x12)) | (~x11 & x12 & x09 & x10)));
  assign z088 = ~x04 & x07 & (x08 ? (x09 & x10 & x11 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & ~x19 & ~x21 & (x01 ? x20 : (~x20 & ~x22))) : (~x09 & ~x10 & (~x11 | ~x12)));
  assign z089 = (x10 & (x09 | x11)) | ~x01 | x04 | ~x07 | x08;
  assign z090 = ~x04 & x07 & x09 & x10 & x11 & ((~x08 & ~x12) | (~x01 & x08 & x12 & ~x13 & ~x14 & ~x15 & ~x16 & ~x17 & x18 & ~x19 & x20 & x21 & x22));
  assign z091 = x21 & x20 & ~x19 & x18 & ~x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & x01 & ~x04;
  assign z092 = x11 & x10 & ~x09 & ~x08 & ~x04 & x07;
  assign z093 = ~x04 & ~x07 & x12 & ((~x08 & ~x09 & x10) | (~x10 & x11 & x08 & x09));
  assign z094 = x23;
  assign z095 = x10 & x09 & ~x08 & ~x04 & ~x07;
  assign z096 = x12 & x11 & x10 & x09 & ~x08 & ~x04 & x07;
  assign z097 = ~x12 & x11 & ~x10 & ~x09 & x08 & ~x04 & x07;
  assign z098 = ~x04 & x07 & x08 & x10 & ((~x11 & x12) | (x09 & x11 & ~x12));
  assign z099 = x12 & x11 & ~x10 & x09 & ~x08 & ~x04 & ~x07;
  assign z100 = ~x04 & ~x07 & x08 & x11 & (~x09 | ~x12);
  assign z101 = x21 & x20 & x19 & ~x18 & x17 & ~x16 & ~x15 & ~x14 & ~x13 & x12 & x11 & x10 & x09 & x08 & x07 & ~x01 & ~x04;
  assign z102 = 1'b0;
  assign z103 = 1'b0;
  assign z104 = 1'b0;
  assign z105 = 1'b0;
  assign z106 = 1'b0;
  assign z107 = 1'b0;
  assign z108 = 1'b0;
endmodule