module pla__t2 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15;
  assign z00 = ~x00 & ~x12 & ((~x14 & ((~x13 & ((x01 & x03 & ~x04 & ~x11 & ~x15 & ~x16 & (x06 | (~x02 & ~x06))) | (x11 & x16))) | (x11 & (~x16 | (x13 & ~x15 & x16))))) | (x11 & ~x13 & x14 & ~x15));
  assign z01 = ~x00 & ~x11 & ((~x13 & (x12 | (x01 & ~x02 & ~x03 & x04 & ~x05 & ~x12 & ~x14 & ~x15 & ~x16))) | (x12 & x13 & (~x14 | (x14 & (~x15 | (x15 & ~x16))))));
  assign z02 = ~x00 & ((x13 & (((~x15 | (x15 & ~x16)) & (x11 ? (~x12 & ~x14) : (x12 & x14))) | (~x11 & x12 & ~x14))) | (~x11 & ~x13 & ((x12 & x14 & x15 & x16) | (x01 & x03 & ~x04 & x06 & ~x15 & ~x16 & ~x12 & ~x14))));
  assign z03 = ~x00 & ((~x12 & ((x11 & ((~x13 & x14 & ~x15) | (~x14 & x15 & x16))) | (~x07 & x10 & ~x11 & ~x15 & ~x16 & ~x13 & x14))) | (~x11 & x12 & (x14 ? (~x15 | (x15 & ~x16)) : (x15 & x16))));
  assign z04 = ~x00 & (x15 ? (~x16 & (x11 ? (~x12 & ~x14) : x12)) : (x16 & (x11 ? (~x12 & (~x13 | (x13 & ~x14))) : ((x12 & (x14 | (x13 & ~x14))) | (~x13 & ~x14)))));
  assign z05 = ~x00 & ~x16 & (x12 ? ~x11 : ((x11 & (~x14 | (~x13 & x14 & ~x15))) | (x01 & ~x03 & x04 & x05 & ~x11 & ~x13 & ~x14 & ~x15)));
  assign z06 = ~x00 & ((~x11 & ((x12 & (((~x15 | (x15 & x16)) & (~x13 | (x13 & x14))) | (x13 & ~x14) | (x14 & x15 & ~x16))) | (~x13 & ~x14 & ~x16 & (x15 | (x01 & ~x12 & ~x15 & (~x02 | (x04 & x05) | (x03 & x06))))))) | (~x12 & ((x11 & ((~x14 & ((x13 & (x16 | (x15 & ~x16))) | (~x15 & ~x16) | (~x13 & x15))) | (~x13 & x14 & (~x15 | (x15 & ~x16))))) | (~x15 & x16 & ~x13 & ~x14))));
  assign z07 = ~x00 & ~x12 & (x11 ? (x13 & ~x14) : (~x13 & ~x15 & ~x16 & (x14 | (x01 & x03 & x06 & ~x14))));
  assign z08 = x07 & ~x11 & ~x12 & ~x13 & ~x14 & (x15 ^ x16);
  assign z09 = (~x13 & ((~x14 & ((~x15 & ((x07 & (x11 ^ x12)) | (~x07 & ~x11 & ~x12 & x16))) | (~x07 & ~x11 & ~x12 & x15 & ~x16))) | (~x07 & x11 & ~x12 & x14 & (x15 ^ x16)))) | (~x07 & ~x11 & x12 & x13 & (x14 ? (~x15 & ~x16) : (x15 & x16)));
  assign z10 = ~x11 & x12 & ((~x13 & x15 & (x16 | (x14 & ~x16))) | (x14 & ~x15) | (x13 & ~x14));
  assign z11 = ~x11 & x12 & ((x13 & (~x14 | (x14 & ~x15 & ~x16))) | (x15 & x16 & ~x13 & x14));
  assign z12 = x07 & x11 & ~x12 & ~x13 & (~x14 ^ ~x15);
  assign z13 = x07 & ~x08 & x11 & ~x12 & ~x13 & (~x14 ^ ~x15);
  assign z14 = x07 & x09 & x11 & ~x12 & ~x13 & (~x14 ^ ~x15);
  assign z15 = x16 & x15 & ~x14 & x13 & ~x12 & x07 & x11;
endmodule