module pla__ts10 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15;
  assign z00 = x16 ? (~x19 & (x17 ? (~x20 & ((x10 & ~x18 & x21) | (x09 & x18 & ~x21))) : (x20 & ((x12 & ~x18 & x21) | (x11 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x14 & ~x18 & x21) | (x13 & x18 & ~x21))) : (x20 & ((x00 & ~x18 & x21) | (x15 & x18 & ~x21)))));
  assign z01 = x16 ? (~x19 & (x17 ? (~x20 & ((x11 & ~x18 & x21) | (x10 & x18 & ~x21))) : (x20 & ((x13 & ~x18 & x21) | (x12 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x15 & ~x18 & x21) | (x14 & x18 & ~x21))) : (x20 & ((x01 & ~x18 & x21) | (x00 & x18 & ~x21)))));
  assign z02 = x16 ? (~x19 & (x17 ? (~x20 & ((x12 & ~x18 & x21) | (x11 & x18 & ~x21))) : (x20 & ((x14 & ~x18 & x21) | (x13 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x00 & ~x18 & x21) | (x15 & x18 & ~x21))) : (x20 & ((x02 & ~x18 & x21) | (x01 & x18 & ~x21)))));
  assign z03 = x16 ? (~x19 & (x17 ? (~x20 & ((x13 & ~x18 & x21) | (x12 & x18 & ~x21))) : (x20 & ((x15 & ~x18 & x21) | (x14 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x01 & ~x18 & x21) | (x00 & x18 & ~x21))) : (x20 & ((x03 & ~x18 & x21) | (x02 & x18 & ~x21)))));
  assign z04 = x16 ? (~x19 & (x17 ? (~x20 & ((x14 & ~x18 & x21) | (x13 & x18 & ~x21))) : (x20 & ((x00 & ~x18 & x21) | (x15 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x02 & ~x18 & x21) | (x01 & x18 & ~x21))) : (x20 & ((x04 & ~x18 & x21) | (x03 & x18 & ~x21)))));
  assign z05 = x16 ? (~x19 & (x17 ? (~x20 & ((x15 & ~x18 & x21) | (x14 & x18 & ~x21))) : (x20 & ((x01 & ~x18 & x21) | (x00 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x03 & ~x18 & x21) | (x02 & x18 & ~x21))) : (x20 & ((x05 & ~x18 & x21) | (x04 & x18 & ~x21)))));
  assign z06 = x16 ? (~x19 & (x17 ? (~x20 & ((x00 & ~x18 & x21) | (x15 & x18 & ~x21))) : (x20 & ((x02 & ~x18 & x21) | (x01 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x04 & ~x18 & x21) | (x03 & x18 & ~x21))) : (x20 & ((x06 & ~x18 & x21) | (x05 & x18 & ~x21)))));
  assign z07 = x16 ? (~x19 & (x17 ? (~x20 & ((x01 & ~x18 & x21) | (x00 & x18 & ~x21))) : (x20 & ((x03 & ~x18 & x21) | (x02 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x05 & ~x18 & x21) | (x04 & x18 & ~x21))) : (x20 & ((x07 & ~x18 & x21) | (x06 & x18 & ~x21)))));
  assign z08 = x16 ? (~x19 & (x17 ? (~x20 & ((x02 & ~x18 & x21) | (x01 & x18 & ~x21))) : (x20 & ((x04 & ~x18 & x21) | (x03 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x06 & ~x18 & x21) | (x05 & x18 & ~x21))) : (x20 & ((x08 & ~x18 & x21) | (x07 & x18 & ~x21)))));
  assign z09 = x16 ? (~x19 & (x17 ? (~x20 & ((x03 & ~x18 & x21) | (x02 & x18 & ~x21))) : (x20 & ((x05 & ~x18 & x21) | (x04 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x07 & ~x18 & x21) | (x06 & x18 & ~x21))) : (x20 & ((x09 & ~x18 & x21) | (x08 & x18 & ~x21)))));
  assign z10 = x16 ? (~x19 & (x17 ? (~x20 & ((x04 & ~x18 & x21) | (x03 & x18 & ~x21))) : (x20 & ((x06 & ~x18 & x21) | (x05 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x08 & ~x18 & x21) | (x07 & x18 & ~x21))) : (x20 & ((x10 & ~x18 & x21) | (x09 & x18 & ~x21)))));
  assign z11 = x16 ? (~x19 & (x17 ? (~x20 & ((x05 & ~x18 & x21) | (x04 & x18 & ~x21))) : (x20 & ((x07 & ~x18 & x21) | (x06 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x09 & ~x18 & x21) | (x08 & x18 & ~x21))) : (x20 & ((x11 & ~x18 & x21) | (x10 & x18 & ~x21)))));
  assign z12 = x16 ? (~x19 & (x17 ? (~x20 & ((x06 & ~x18 & x21) | (x05 & x18 & ~x21))) : (x20 & ((x08 & ~x18 & x21) | (x07 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x10 & ~x18 & x21) | (x09 & x18 & ~x21))) : (x20 & ((x12 & ~x18 & x21) | (x11 & x18 & ~x21)))));
  assign z13 = x16 ? (~x19 & (x17 ? (~x20 & ((x07 & ~x18 & x21) | (x06 & x18 & ~x21))) : (x20 & ((x09 & ~x18 & x21) | (x08 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x11 & ~x18 & x21) | (x10 & x18 & ~x21))) : (x20 & ((x13 & ~x18 & x21) | (x12 & x18 & ~x21)))));
  assign z14 = x16 ? (~x19 & (x17 ? (~x20 & ((x08 & ~x18 & x21) | (x07 & x18 & ~x21))) : (x20 & ((x10 & ~x18 & x21) | (x09 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x12 & ~x18 & x21) | (x11 & x18 & ~x21))) : (x20 & ((x14 & ~x18 & x21) | (x13 & x18 & ~x21)))));
  assign z15 = x16 ? (~x19 & (x17 ? (~x20 & ((x09 & ~x18 & x21) | (x08 & x18 & ~x21))) : (x20 & ((x11 & ~x18 & x21) | (x10 & x18 & ~x21))))) : (x19 & (x17 ? (~x20 & ((x13 & ~x18 & x21) | (x12 & x18 & ~x21))) : (x20 & ((x15 & ~x18 & x21) | (x14 & x18 & ~x21)))));
endmodule