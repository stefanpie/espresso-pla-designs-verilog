module pla__apex3 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49;
  assign z00 = (~x48 & ((x50 & ((~x53 & ((x49 & ((x11 & ((x46 & ~x47 & ~x51 & x52) | (~x46 & x47 & ~x52))) | (x46 & ~x47 & (x51 ? x52 : (~x52 | (x52 & (x10 | x25 | (~x10 & ~x11 & ~x25)))))))) | (~x49 & (x46 ? (~x47 & (~x21 | (x21 & x51 & x52))) : (x47 & ((x51 & x52) | (x28 & ~x51 & ~x52))))) | (x46 & ~x47 & x51 & ~x52))) | (x49 & ((~x46 & x47 & (x51 ? (x52 & x53) : ~x52)) | (x06 & x46 & ~x47 & x51 & ~x52 & x53))) | (x46 & ~x47 & ((x51 & x52 & x53) | (~x49 & ((x53 & (~x51 | (~x22 & ~x25 & ~x28 & x51 & ~x52))) | (x51 & ~x52 & (x22 | x25 | x28)))))))) | (~x50 & ((~x47 & ((~x51 & ((~x49 & x52 & x53) | (x46 & x49 & ~x53))) | (x46 & (x49 ? (x51 & (x52 | (~x52 & (x24 | ~x53 | (~x24 & x53))))) : ((~x52 & x53) | (~x39 & x51 & x52)))) | (~x46 & x49 & x51 & x53))) | (~x46 & ((x47 & ((~x53 & (x52 ? (x51 | (x31 & ~x49 & ~x51)) : ((x49 & (~x51 | (~x20 & x51))) | (x09 & ~x51) | (~x49 & x51)))) | (x39 & ~x49 & ~x51 & ~x52 & x53))) | (x13 & ~x49 & ~x51 & x52 & x53))))) | (x46 & ~x47 & ~x51 & (~x49 ^ x53)))) | (x48 & ((~x47 & ((~x49 & ((x46 & ((~x53 & (x50 ? (x52 & (x51 ? ~x03 : ~x04)) : ((~x52 & ((~x37 & x51 & (x38 | x43)) | (x20 & ~x51))) | (~x16 & ~x51 & x52)))) | (~x04 & ((x50 & ~x51 & ~x52) | (x52 & x53 & ~x50 & x51))) | (x50 & x52 & x53))) | (x40 & ~x46 & ~x50 & x51 & ~x52 & ~x53))) | (~x46 & x49 & x51 & ((x50 & ~x52 & (x53 ? x41 : x07)) | (~x34 & ~x50 & x52 & ~x53))))) | (~x46 & x47 & x52 & ((x49 & (x53 ? x51 : x50)) | (~x49 & x50 & ~x51 & x53))))) | (~x47 & ~x50 & x51 & x52 & ((x49 & x53 & x17 & ~x46) | (x46 & ~x49 & ~x53)));
  assign z01 = x46 ? (~x47 & ~x49 & ((x51 & ((~x50 & ((~x48 & ((~x52 & ~x53) | (x39 & x52 & x53))) | (~x52 & ~x53 & (x37 | (~x38 & ~x43))) | (x52 & x53 & x04 & x48))) | (x48 & ((~x52 & x53) | (x50 & ~x53 & (~x52 | (x03 & x52))))))) | (x48 & ~x51 & ((x04 & x50 & (~x52 | (x52 & ~x53))) | (~x50 & (x53 | (x16 & x52 & ~x53))))))) : ((x53 & ((x29 & ((x47 & ~x48 & ~x49 & ~x50 & x51) | (x50 & ~x51 & ~x52 & ~x47 & x48 & x49))) | (x47 & ((~x51 & ((~x38 & ((~x48 & x49 & ~x50 & x52) | (x01 & x43 & x48 & ~x52))) | (x49 & (~x50 ^ x52)) | (x48 & ((~x50 & x52) | (~x49 & ~x52 & (x50 | (~x50 & (~x01 | x38 | ~x43)))))) | (~x50 & ~x52 & ~x39 & ~x48))) | (~x48 & ((x51 & ((x49 & (~x50 | (x50 & ~x52))) | (~x29 & ~x50 & ~x52) | (~x49 & x52))) | (~x49 & x50 & ~x52))) | (~x50 & x52 & ~x13 & ~x49) | (x48 & x49 & ~x52))) | (~x47 & ((x48 & x51 & (x49 ? (x50 & x52) : (~x50 & ~x52))) | (x41 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52))))) | (x47 & ((~x53 & (x48 ? ((~x50 & ((x01 & (x49 ? x51 : (~x51 & ~x52))) | (x49 & (~x51 | (x51 & (~x43 | x52)))))) | (~x51 & ((x50 & ~x52) | (~x49 & (~x01 | x52)))) | (x51 & ~x52 & x49 & x50)) : ((x50 & ((x51 & (x49 ? (x52 | (~x11 & ~x52)) : ~x52)) | (~x28 & ~x49 & ~x51))) | (~x51 & ((x52 & (~x31 | x49)) | (~x50 & ~x52 & ~x09 & ~x49)))))) | (x51 & ((x48 & (~x49 | (x49 & ~x52 & ~x01 & x43))) | (~x50 & ~x52 & x20 & x49))) | (~x48 & ~x51 & x52 & ((~x49 & x50) | (x38 & x49 & ~x50))))) | (~x47 & x48 & x51 & x52 & ~x53 & ((x39 & x49 & x50) | (~x49 & ~x50))));
  assign z02 = x48 ? ((~x47 & ((~x49 & (x46 ? ((~x04 & ((x50 & ~x51 & ~x52) | (x52 & x53 & ~x50 & x51))) | (x51 & ((x50 & x52 & x53) | (~x53 & ((~x52 & (x50 | (~x37 & ~x50 & (x38 | x43)))) | (~x03 & x50 & x52))))) | (~x51 & ((x52 & ~x53) | (~x52 & x53 & x04 & x50)))) : ((x52 & ((~x50 & (~x51 ^ x53)) | (x20 & x51 & x53))) | (~x50 & ~x51 & (x53 | (x37 & ~x52 & ~x53)))))) | (~x46 & x49 & (x52 ? ((~x51 & ((~x50 & (~x20 | (x20 & ~x53))) | x53 | (~x29 & x50))) | (x51 & ((x50 & (~x53 | (x42 & x53))) | (~x17 & ~x50 & x53))) | (x29 & x50 & ~x53)) : (~x53 | (x51 & x53 & x19 & ~x50)))))) | (~x46 & ((x47 & ((~x52 & ((~x51 & ((x01 & ((~x38 & x43 & x53) | (~x49 & ~x50 & ~x53))) | (x50 & (x49 | ~x53)) | (~x49 & ~x50 & x53 & (~x01 | x38 | ~x43)))) | (x49 & x51 & ((~x01 & x43) | x53 | (x50 & ~x53))))) | (~x51 & ((x49 & (x50 ? (x52 & x53) : ~x53)) | (x52 & (x53 ? ~x50 : ~x49)) | (~x49 & (x53 ? x50 : ~x01)))) | (x51 & (~x49 | (x49 & ~x50 & (x52 | (~x53 & (x01 | ~x43)))))))) | (x50 & ((~x49 & ((~x52 & x53 & x29 & ~x51) | (x51 & x52 & ~x53))) | (~x52 & ((x51 & x53 & ~x41 & x49) | (x08 & ~x51 & ~x53))))) | (x49 & ~x51 & ~x52 & x53 & (~x29 | ~x50))))) : ((x49 & ((~x47 & ((~x51 & (x46 ? (x50 ? (~x52 & x53) : (x52 & ~x53)) : (x50 & x52 & (x53 ? x20 : x08)))) | (x50 & x51 & ((x52 & ((x03 & x53) | (x30 & ~x46 & ~x53))) | (~x46 & ~x52 & (x53 ? x44 : x35)))))) | (~x46 & x47 & ((~x52 & (x50 ? (x53 & (~x51 | (~x43 & x51))) : (~x53 & (~x51 | (~x20 & x51))))) | (x50 & x52 & x53 & (x51 | (~x01 & ~x51))))))) | (~x49 & ((~x47 & ~x50 & ((x46 & x51 & ((~x52 & ~x53) | (x39 & x52 & x53))) | (~x52 & x53 & ~x46 & ~x51))) | (x28 & ~x46 & x47 & ~x52 & ~x53 & x50 & ~x51))) | (x51 & x52 & ~x53 & ~x46 & x47 & ~x50));
  assign z03 = (~x46 & ((x51 & ((x48 & ((~x52 & ((x47 & ((~x01 & (x49 ? x43 : (x50 & ~x53))) | (x50 & (x53 ? x43 : (x49 | (~x26 & ~x49)))))) | (x50 & ((~x47 & (~x49 | (~x07 & x49 & ~x53))) | (~x41 & x49 & x53))) | (~x47 & ~x50 & (x53 | (~x40 & ~x49 & ~x53))))) | (x49 & ((x52 & (x47 ? ~x53 : (x50 ? (~x53 | (x42 & x53)) : (x53 ? ~x17 : ~x34)))) | (x47 & ~x50 & ~x53 & (x01 | ~x43)))) | (x50 & x52 & x53 & x45 & x47 & ~x49))) | (~x48 & (x50 ? (x49 ? (~x52 & ((x47 & (x53 ? x43 : ~x11)) | (~x35 & ~x53) | (~x44 & ~x47 & x53))) : (x47 ? x52 : ((~x14 & x53) | (~x16 & x52 & ~x53)))) : ((x49 & (x53 | (~x47 & ~x52 & (~x41 | (x41 & ~x53))))) | (~x52 & ~x53 & x47 & ~x49)))) | (x52 & ((~x47 & x53 & ((~x49 & x50) | (x17 & x49 & ~x50))) | (x50 & ~x53 & ~x30 & x49))) | (x20 & x47 & x49 & ~x50 & ~x52))) | (~x51 & ((x47 & ((x01 & ((x50 & x52 & x53 & ~x48 & x49) | (x48 & ~x49 & ~x50 & ~x52 & ~x53))) | (x49 & ~x50 & ((~x48 & x52 & (x38 | (~x38 & x53))) | (~x52 & x53) | (x48 & ~x53))))) | (~x53 & (x50 ? ((~x08 & (x48 ? ~x47 : (x49 & x52))) | (x49 & ~x52) | (x48 & x52)) : ((~x48 & x49 & x52) | (~x47 & (x48 ? ((x20 & x49 & x52) | (~x37 & ~x49 & ~x52)) : (x49 & ~x52)))))) | (~x47 & ((x49 & ((x52 & ((~x20 & (x50 ? x53 : x48)) | (x48 & x53))) | (~x52 & x53 & ~x48 & x50))) | (x53 & ((~x48 & ~x49 & ~x50 & (x52 | (x41 & ~x52))) | (~x29 & x48 & x50))))) | (x48 & x49 & ~x50 & ~x52 & x53))) | (x49 & ((x47 & (x48 ? (x53 & (~x52 | (x50 & x52))) : (x50 & ~x53 & (x52 | (x11 & ~x52))))) | (~x50 & ~x52 & ~x53 & ~x47 & x48))))) | (~x47 & ((x46 & ((~x49 & ((x48 & ((x04 & ((x52 & x53 & ~x50 & x51) | (x50 & ~x51 & ~x53))) | (~x50 & ~x51 & (x52 ? (x53 | (x16 & ~x53)) : ~x53)) | (x51 & x52 & ~x53 & x03 & x50))) | (~x48 & ((x53 & (x50 ? x52 : ((~x51 & ~x52) | (x39 & x51 & x52)))) | (x51 & ~x52 & ~x53) | (x50 & ((x51 & ~x52 & (x22 | x25 | x28)) | (~x53 & (~x21 | ~x51)))))) | (~x50 & x51 & ~x52 & ~x53 & (x37 | (~x38 & ~x43))))) | (~x48 & x49 & ((x53 & ((~x51 & x52) | (x51 & ~x52 & ~x24 & ~x50))) | (x51 & (x50 ? (~x52 | (x52 & ~x53)) : (x52 | (~x52 & (x24 | ~x53))))) | (~x51 & ~x53 & (~x52 | (x50 & x52 & (x25 | (~x10 & ~x11 & ~x25) | x10 | x11)))))))) | (x52 & ((x48 & ~x49 & (x50 ? (~x51 & x53) : (x51 & ~x53))) | (~x03 & ~x48 & x49 & x50 & x51 & x53))) | (~x51 & ~x52 & x53 & ~x48 & x49 & ~x50)));
  assign z04 = (x50 & ((~x46 & ((x47 & ((x01 & ((~x51 & x52 & x53 & ~x48 & x49) | (x51 & ~x53 & x26 & ~x49))) | (~x48 & (x49 ? ((~x52 & ((x51 & (x53 ? x43 : ~x11)) | (x11 & ~x53))) | (~x51 & x52 & ~x53)) : (x53 ? ~x52 : (x52 | (~x28 & ~x51))))) | (x48 & ((x49 & (~x51 | (x51 & ~x53))) | (~x49 & ((~x51 & ~x52 & x53) | (~x45 & x51 & x52))) | (~x52 & ((~x51 & ~x53) | (~x43 & x51 & x53))))) | (x52 & x53 & ~x49 & ~x51))) | (~x53 & ((~x51 & ((~x08 & (x48 ? ~x47 : (x49 & x52))) | (~x52 & (x49 | (x08 & x48))))) | (x51 & (x49 ? ((~x47 & (x48 ? (x52 | (~x07 & ~x52)) : (x52 ? x30 : x35))) | (~x30 & x52) | (~x35 & ~x48 & ~x52)) : (x48 ? x52 : (~x52 | (x16 & ~x47 & x52))))) | (x29 & ~x47 & x48 & x49 & x52))) | (~x47 & ((~x20 & ((x48 & ~x49) | (x52 & x53 & x49 & ~x51))) | (x48 & ((~x51 & ((~x29 & (x53 | (x49 & x52))) | (x52 & (~x49 | (x49 & x53))))) | (x49 & x51 & x53 & (x52 ? x42 : x41)))) | (~x48 & x53 & (x49 ? (~x52 | (x20 & ~x51 & x52)) : ~x51)))) | (~x52 & ((x48 & x53 & ((~x41 & x49 & x51) | (x29 & ~x49 & ~x51))) | (~x49 & x51 & x14 & ~x48))))) | (~x47 & (x51 ? (x52 ? ((~x03 & ((~x48 & x49 & x53) | (~x49 & ~x53 & x46 & x48))) | (x46 & (x48 ? (~x49 & x53) : (~x53 & (x49 | (x21 & ~x49)))))) : ((x48 & ~x49) | (x46 & ~x48 & (x49 | ~x53 | (~x49 & (x22 | x25 | x28 | (~x22 & ~x25 & ~x28 & x53))))))) : ((x46 & ((~x49 & (x48 ? (x52 ? ~x53 : ~x04) : (x53 & (x52 | (x41 & ~x52))))) | (~x48 & x49 & (x53 | (~x53 & (~x52 | (x52 & (x25 | (~x10 & ~x11 & ~x25) | x10 | x11)))))))) | (~x48 & ~x49 & ~x53)))))) | (~x50 & ((~x47 & ((~x49 & ((x52 & ((x16 & ((x51 & x53 & ~x46 & ~x48) | (~x51 & ~x53 & x46 & x48))) | (x51 & ((x46 & ~x48 & (~x39 | (x39 & x53))) | (x48 & x53 & x03 & ~x46))))) | (x46 & ((~x48 & (x51 ? ~x53 : (~x52 & x53))) | (~x52 & (x51 ? (~x53 & (x37 | (~x38 & ~x43))) : x48)))) | (~x46 & x48 & ((x51 & (~x53 | (~x52 & x53))) | (~x52 & ~x53 & ~x37 & ~x51))))) | (x49 & x51 & ((~x48 & (x52 ? x53 : (x46 ? (x24 | ~x53) : x53))) | (~x46 & ((x48 & ((x52 & (x53 ? ~x17 : ~x34)) | (~x19 & ~x52 & x53))) | (x17 & x52 & x53))))) | (~x51 & x52 & x53 & ~x46 & ~x48))) | (~x46 & ((~x49 & ((x52 & ((~x48 & ~x51 & ((x13 & x53) | (x31 & x47 & ~x53))) | (x47 & x51 & (~x27 | x53)))) | (x29 & x47 & ~x48 & x51 & x53))) | (x47 & x51 & ((~x21 & x48 & x53) | (~x20 & ~x48 & x49 & ~x52 & ~x53))))))) | (x48 & x53 & ((x49 & x51 & ~x46 & x47) | (x46 & ~x47 & ~x49 & ~x51 & x52))) | (~x46 & x47 & ~x48 & x51 & ((x49 & x52) | (~x52 & ~x53 & ~x31 & ~x49)));
  assign z05 = (~x47 & ((x51 & ((x53 & ((x52 & ((~x03 & ((~x48 & x49 & x50) | (~x49 & ~x50 & ~x46 & x48))) | (x48 & ((x46 & ~x49 & (x50 | (~x04 & ~x50))) | (x49 & x50 & x42 & ~x46))) | (~x46 & ~x50 & ((~x48 & (x49 | (~x16 & ~x49))) | (x17 & x49))))) | (~x52 & ((~x48 & (x46 ? ((x49 & (x50 ? x06 : ~x24)) | (~x22 & ~x25 & ~x28 & ~x49 & x50)) : (~x49 | (x49 & x50)))) | (x19 & ~x46 & x48 & x49 & ~x50))) | (~x14 & ~x46 & ~x48 & ~x49 & x50))) | (~x53 & ((~x49 & (x46 ? ((x48 & (x50 | (~x37 & ~x50 & ~x52 & (x38 | x43)))) | (x50 & x52 & x21 & ~x48)) : (~x48 & (~x50 | (x50 & (~x52 | (x16 & x52))))))) | (~x48 & (x46 ? (~x52 | (x49 & x52)) : (x49 & ((x30 & x50 & x52) | (x41 & ~x50 & ~x52))))) | (~x46 & x48 & x49 & x52 & (x50 ? ~x39 : ~x34)))) | (~x48 & ~x52 & ((x49 & ~x50 & (x46 ? x24 : ~x41)) | (x46 & ~x49 & x50 & (x22 | x25 | x28)))))) | (~x51 & ((x20 & ((x50 & x52 & x53 & ~x46 & ~x48 & x49) | (~x50 & ~x52 & ~x53 & x46 & x48 & ~x49))) | (x52 & ((x49 & (x46 ? (~x48 & (~x50 | (x50 & ~x53 & (x10 | x11 | x25)))) : ((~x20 & (x50 ? x53 : x48)) | (x50 & ((x48 & (~x29 | x53)) | (x08 & ~x48 & ~x53)))))) | (~x50 & ((~x46 & (x53 | (~x49 & ~x53 & x32 & ~x48))) | (~x49 & ((~x48 & x53) | (x48 & ~x53 & x16 & x46))))) | (x46 & ~x48 & ~x49 & (~x36 | (x50 & x53))))) | (~x52 & ((x50 & (x46 ? (~x49 & ((x04 & x48) | (~x41 & ~x48 & x53))) : (x49 & x53 & (x48 ? x29 : x37)))) | (~x46 & ~x48 & ~x50 & x53 & (~x49 | (~x14 & x49))))) | (~x49 & x50 & ~x53 & x46 & ~x48))) | (~x50 & ((~x52 & x53 & x46 & ~x49) | (~x46 & ~x48 & x49 & x52 & ~x53))))) | (~x46 & ((x47 & ((x48 & ((x53 & ((~x52 & ((~x43 & ((x50 & x51) | (~x49 & ~x50 & ~x51))) | (~x49 & ~x50 & (x51 ? x21 : (~x01 | x38))))) | (x50 & (x51 ? x49 : x52)) | (~x49 & ~x50 & x52))) | (x52 & ((~x53 & ((x49 & (x50 | (~x50 & x51))) | (x27 & ~x50 & x51))) | (x50 & x51 & ~x45 & ~x49))) | (x01 & ~x49 & ~x50 & ~x51 & ~x52 & ~x53))) | (x50 & ((x01 & ((~x51 & x52 & x53 & ~x48 & x49) | (x51 & ~x53 & x26 & ~x49))) | (~x48 & ((x51 & (x53 ? ~x52 : (~x49 | (x49 & (x52 | (~x11 & ~x52)))))) | (~x52 & ~x53 & x11 & x49))))) | (~x48 & ((~x51 & ((x49 & ((~x52 & ~x53) | (x52 & x53 & ~x38 & ~x50))) | (x31 & ~x49 & ~x50 & x52 & ~x53))) | (~x50 & x51 & ((~x49 & x52) | (~x29 & ~x52 & x53))))) | (~x50 & ((x51 & ~x52 & ~x53) | (x52 & x53 & ~x13 & ~x49))))) | (~x48 & (x49 ? (x51 & ~x52 & ((~x50 & x53) | (~x35 & x50 & ~x53))) : (~x51 & x52 & x53 & (x50 | (x13 & ~x50))))) | (x51 & ((x48 & x50 & (x49 ? (~x52 & (~x53 | (~x41 & x53))) : (x52 & ~x53))) | (~x50 & ~x52 & ~x53 & x12 & x49)))));
  assign z06 = (~x46 & ((~x52 & ((x53 & ((x47 & ((x48 & ((x01 & (x49 | (~x38 & x43 & ~x51))) | (~x49 & ((x50 & ~x51) | (x21 & ~x50 & x51))) | (x49 & ~x51) | (~x43 & x50 & x51))) | (~x48 & ((x51 & ((x49 & (~x50 | (x43 & x50))) | (~x29 & ~x50))) | (~x49 & (x50 | (x39 & ~x50 & ~x51))) | (~x39 & ~x50 & ~x51))) | (x49 & ~x50 & ~x51))) | (x49 & ((~x47 & ((~x48 & ((~x44 & x50 & x51) | (~x14 & ~x50 & ~x51))) | (~x50 & x51 & x19 & x48))) | (x50 & ((~x41 & x48 & x51) | (~x48 & ~x51))) | (x48 & ~x51 & (~x29 | ~x50)))) | (~x49 & ((~x47 & ~x50 & (~x51 | (x48 & x51))) | (x50 & ~x51 & x29 & x48))))) | (x51 & (x47 ? ((x48 & ((~x01 & (x49 ? x43 : (x50 & ~x53))) | (x50 & ~x53 & (x49 | (~x26 & ~x49))))) | (~x20 & ~x48 & x49 & ~x50 & ~x53)) : (~x53 & ((~x48 & ((x49 & (x50 ? x35 : x41)) | (x25 & ~x49 & x50))) | (~x49 & ~x50 & x40 & x48))))) | (~x48 & x49 & ~x50 & ~x51 & ~x53 & (x47 | (x25 & ~x47))))) | (~x48 & ((~x14 & ((x50 & x51 & x53 & ~x47 & ~x49) | (x52 & ~x53 & x49 & ~x51))) | (x52 & ((~x53 & ((x25 & ((x50 & ~x51) | (~x47 & ~x49 & x51))) | (~x47 & ((~x49 & ((x50 & x51) | (~x32 & ~x50 & ~x51))) | (x50 & ~x51 & x08 & x49))) | (x50 & ((x47 & (~x51 | (x49 & x51))) | (~x08 & x49 & ~x51))) | (~x31 & x47 & ~x51))) | (x49 & ~x51 & ((x38 & x47 & ~x50) | (x50 & x53 & x20 & ~x47))))))) | (x48 & ((~x47 & ((x52 & ((~x50 & ((~x53 & (x49 ? (x51 ? x34 : x20) : ~x51)) | (x51 & x53 & ~x03 & ~x49))) | (x49 & x50 & ((x29 & ~x53) | (x51 & (~x53 | (x42 & x53))))))) | (~x15 & x49 & ~x50 & ~x51 & x53))) | (x52 & ((x47 & ((x51 & ((~x49 & x50 & (~x45 | (x45 & x53))) | (~x50 & (x49 | (x27 & ~x53))))) | (~x49 & ~x51 & ~x53))) | (~x49 & x50 & x51 & ~x53))))) | (~x51 & x52 & ~x53 & x47 & x49 & ~x50))) | (~x47 & ((x51 & (x52 ? ((x50 & ((~x03 & ((~x48 & x49 & x53) | (~x49 & ~x53 & x46 & x48))) | (x46 & ~x48 & ~x53 & (x49 | (x21 & ~x49))))) | (x46 & ~x49 & ~x50 & (~x53 | (x53 & (x48 ? ~x04 : x39))))) : ((x46 & ((~x48 & ((~x49 & ~x50 & ~x53) | (x53 & ((x49 & (x50 ? x06 : ~x24)) | (~x22 & ~x25 & ~x28 & ~x49 & x50))))) | (~x49 & ((x48 & x53) | (~x50 & ~x53 & (x37 | (~x38 & ~x43))))))) | (~x48 & ~x49 & ~x50 & x53)))) | (x46 & ((~x51 & (x48 ? (~x49 & ~x53 & (x50 ? (x04 ^ x52) : (x52 ? ~x16 : x20))) : ((x49 & (x50 ? ((~x52 & x53) | (~x10 & ~x11 & ~x25 & x52 & ~x53)) : ~x52)) | (x14 & ~x49 & ~x50 & x52 & x53)))) | (x52 & ((~x48 & ~x50 & ~x53 & (x36 | x49)) | (x50 & x53 & x48 & ~x49))))) | (~x51 & ~x52 & x53 & ~x48 & ~x49 & x50)));
  assign z07 = (~x46 & ((~x53 & ((x47 & ((x51 & ((x01 & ((x48 & x49 & ~x50) | (x26 & ~x49 & x50))) | (x48 & ((~x50 & ((x49 & (~x43 | x52)) | (x27 & x52))) | (~x49 & x50 & ~x52 & (~x01 | ~x26)))) | (~x48 & (x49 ? ((x50 & (x52 | (~x11 & ~x52))) | (~x20 & ~x50 & ~x52)) : (x50 ^ x52))) | (~x49 & (x52 ? x50 : x05)))) | (~x51 & ((x49 & (~x48 | (x48 & ~x50 & ~x52))) | (~x49 & (x48 ? (~x01 | x52) : ((~x52 & (x50 ? x28 : ~x09)) | (x50 & (~x28 | x52))))) | (x48 & (x52 ? x05 : x50)) | (~x31 & ~x48 & x52))) | (x49 & x50 & ((x48 & x52) | (x11 & ~x48 & ~x52))))) | (x50 & ((~x51 & ((x08 & ((x48 & ~x52) | (x49 & x52 & ~x47 & ~x48))) | (~x48 & ((~x47 & ~x49) | (~x08 & x49 & x52))) | (x18 & x49 & ~x52))) | (x29 & ~x47 & x48 & x49 & x52) | (x51 & ((~x47 & ((x49 & (x48 ? (x52 | (~x07 & ~x52)) : (x52 ? x30 : x35))) | (~x48 & ~x49 & (x52 | (~x25 & ~x52))))) | (x03 & x48 & x52) | (x49 & ~x52 & ~x35 & ~x48))))) | (x49 & ((~x51 & ((~x47 & ((x48 & (~x52 | (x20 & ~x50 & x52))) | (~x50 & ~x52 & ~x25 & ~x48))) | (~x14 & ~x48 & x52))) | (~x47 & x48 & ~x50 & x51 & (~x52 | (~x34 & x52))))) | (~x50 & ((~x47 & ((x52 & (x48 ? ~x49 : (x51 | (~x32 & ~x49 & ~x51)))) | (x48 & ~x49 & ~x52 & (x51 ? x40 : x37)))) | (x51 & ~x52 & ~x48 & ~x49))))) | (x53 & ((~x47 & ((~x48 & ((~x14 & ((~x49 & x50 & x51) | (~x51 & ~x52 & x49 & ~x50))) | (x49 & ((~x50 & x51) | (~x51 & ~x52 & x37 & x50))) | (~x50 & x52 & (~x51 | (~x16 & ~x49 & x51))))) | (x48 & ((x51 & ((~x50 & ((~x49 & (~x52 | (~x03 & x52))) | (x19 & x49 & ~x52))) | (x49 & x50 & (x52 ? x42 : x41)))) | (x50 & ~x51 & ~x52 & x29 & x49))) | (x17 & x49 & ~x50 & x51 & x52))) | (x47 & ((~x52 & ((~x43 & ((~x48 & x49 & x50 & x51) | (x48 & ~x49 & ~x50 & ~x51))) | (x48 & ~x49 & ~x50 & ~x51 & (~x01 | x38)))) | (x50 & x51 & x52 & (x49 | (x45 & x48 & ~x49))))) | (x13 & ~x48 & ~x49 & ~x50 & ~x51 & x52))) | (x47 & ((x50 & ((~x49 & ((~x52 & ((x43 & (~x48 ^ ~x51)) | (~x51 & (x48 ? ~x26 : (~x00 | ~x23))))) | (x51 & x52 & ~x45 & x48))) | (x49 & x52 & x02 & x48))) | (~x50 & ~x51 & x52 & x38 & ~x48 & x49))) | (~x41 & ~x47 & ~x48 & x51 & ~x52 & x49 & ~x50))) | (~x47 & ((x46 & ((~x49 & ((x50 & ((~x53 & (x48 ? ((x03 & x51 & x52) | (x04 & ~x51 & ~x52)) : (~x21 | (x21 & x51 & x52)))) | (~x48 & ((~x51 & x53 & (x52 | (x41 & ~x52))) | (x51 & ~x52 & (x22 | x25 | x28)) | (x27 & x52))))) | (x48 & ((~x51 & ~x52 & x53) | (~x50 & x52))) | (~x50 & x53 & ((x51 & (~x52 | (x39 & ~x48 & x52))) | (~x48 & ~x51 & (~x52 | (x14 & x52))))) | (~x48 & ~x51 & ~x53))) | (~x48 & ((x49 & (x51 ? (~x53 & (~x20 | ~x50)) : ((~x52 & ~x53) | (x50 & ((~x52 & x53) | (~x10 & ~x11 & ~x25 & x52 & ~x53)))))) | (~x52 & ~x53 & x50 & x51))))) | (~x49 & ((x48 & ~x50 & ((~x29 & ~x52 & x53) | (x26 & ~x51 & x52))) | (~x51 & ~x52 & ~x53 & ~x33 & ~x48))) | (~x03 & ~x48 & x49 & x52 & x53 & x50 & x51)));
  assign z08 = (~x47 & ((x50 & ((~x52 & ((~x48 & ((x46 & ((x51 & ~x53) | (~x49 & ~x51 & x53))) | (~x46 & x49 & ~x51 & x53))) | (~x46 & x48 & ~x49 & x51 & ~x53))) | (~x51 & x52 & x53 & ~x46 & x48 & ~x49))) | (~x46 & ~x49 & ~x50 & ((~x52 & x53 & x48 & x51) | (x52 & ~x53 & ~x48 & ~x51))))) | (~x46 & x47 & ~x48 & x52 & ~x53 & (x49 ? (x50 & ~x51) : (~x50 & x51)));
  assign z09 = ~x46 & ~x51 & x53 & ((x49 & x50 & x52 & x47 & x48) | (~x49 & ~x50 & ~x52 & ~x47 & ~x48));
  assign z10 = ~x46 & ~x49 & ((~x47 & ((~x50 & x51 & (x48 ? (x52 ^ x53) : (~x52 & ~x53))) | (~x51 & x52 & x53 & ~x48 & x50))) | (x51 & x52 & ~x53 & x47 & ~x48 & ~x50));
  assign z11 = (~x46 & x47 & ~x48 & x52 & ~x53 & (x49 ? (x50 & ~x51) : (~x50 & x51))) | (~x47 & ((x51 & ((~x48 & (x46 ? ((x52 & x53 & x49 & ~x50) | (~x52 & ~x53 & ~x49 & x50)) : (~x49 & ~x53 & (~x50 ^ x52)))) | (~x46 & x48 & ~x49 & ~x50 & (x52 ^ x53)))) | (~x46 & ~x48 & ~x49 & x52 & x53 & x50 & ~x51)));
  assign z12 = ~x46 & x47 & ((x53 & ((x51 & ((~x48 & x50 & (~x52 | (x49 & x52))) | (x48 & x49 & ~x50 & x52))) | (x48 & ~x51 & (x49 ? ~x52 : (~x50 & x52))))) | (~x48 & x49 & ~x53 & (x52 ? ~x50 : ~x51)));
  assign z13 = x53 & x52 & ~x51 & ~x50 & ~x49 & ~x48 & ~x46 & ~x47;
  assign z14 = ~x53 & ~x52 & ~x51 & x50 & x49 & x48 & ~x46 & ~x47;
  assign z15 = x50 ? ((~x47 & ((x46 & ~x49 & ((~x51 & x52 & ~x53) | (x48 & (x51 ? (x52 & ~x53) : ~x52)))) | (x51 & x52 & x53 & ~x48 & x49))) | (x51 & x52 & ~x53 & ~x46 & x48 & ~x49)) : ((~x46 & ((x47 & ((x52 & ~x53 & x49 & ~x51) | (x51 & ~x52 & x48 & ~x49))) | (~x51 & ~x52 & ~x53 & ~x47 & x48 & ~x49))) | (~x47 & x48 & ~x49 & x53 & ((x51 & x52) | (x46 & ~x51 & ~x52))));
  assign z16 = (~x48 & ((~x49 & x52 & ((~x47 & ((x46 & (x50 ? (~x51 & x53) : (x51 & ~x53))) | (~x46 & ~x50 & ~x51 & x53))) | (~x46 & x47 & x50 & x51 & ~x53))) | (~x46 & x47 & x49 & x50 & ~x52 & ((x51 & (x53 | (~x11 & ~x53))) | (~x53 & (x11 | ~x51)))))) | (x48 & x49 & ~x46 & x47 & x52 & ~x53 & x50 & ~x51);
  assign z17 = ~x47 & ~x49 & x52 & ((~x46 & ~x48 & x51 & (~x50 ^ ~x53)) | (x46 & x48 & ~x50 & ~x51 & ~x53));
  assign z18 = x46 ? (~x47 & ((~x51 & ~x52 & x53 & ~x48 & x49 & ~x50) | (~x49 & x51 & ((x48 & ~x53 & (x50 ^ x52)) | (x52 & x53 & ~x48 & x50))))) : (x47 & ~x49 & x50 & ~x53 & ((~x48 & (x51 ^ x52)) | (~x51 & ~x52 & x23 & x48)));
  assign z19 = x46 ? (~x47 & ~x48 & x49 & ~x53 & (x50 ? (~x51 & x52 & (x25 | (~x10 & ~x11 & ~x25) | x10 | x11)) : (x51 & ~x52))) : ((~x49 & (x47 ? ((x48 & x53 & (x50 ? (~x51 & ~x52) : (x51 & x52))) | (x51 & ~x52 & ~x53 & ~x48 & x50)) : (~x48 & ((x50 & (x51 ? (~x52 & x53) : (x52 & ~x53))) | (~x50 & x51 & x52 & ~x53))))) | (~x47 & ~x48 & x49 & ~x52 & x53 & ~x50 & ~x51));
  assign z20 = ~x46 & ~x47 & x48 & x49 & ~x50 & x51 & (x52 ^ x53);
  assign z21 = x51 & ((x46 & ~x47 & ~x48 & ~x52 & x53 & ~x49 & ~x50) | (~x46 & x47 & x48 & x52 & ~x53 & x49 & x50));
  assign z22 = (~x46 & ((x49 & ((~x51 & ((x47 & x52 & x53 & (~x48 ^ ~x50)) | (~x50 & ~x52 & ~x53 & ~x47 & ~x48))) | (x51 & ~x52 & x53 & ~x47 & x48 & ~x50))) | (~x52 & ~x53 & x50 & x51 & ~x47 & ~x48 & ~x49))) | (~x52 & ~x53 & x50 & ~x51 & x46 & ~x47 & ~x48 & x49);
  assign z23 = ~x53 & x52 & x51 & x50 & ~x49 & ~x46 & x47;
  assign z24 = ~x48 & x49 & x52 & ~x53 & ((x46 & ~x47 & ~x50 & x51) | (~x46 & x47 & x50 & ~x51));
  assign z25 = ~x46 & ~x47 & x48 & x49 & ~x50 & (x51 ? ~x52 : (x52 & x53));
  assign z26 = ~x51 & x52 & ((~x46 & x47 & ~x49 & x50 & x53) | (x49 & ~x50 & ~x53 & x46 & ~x47 & ~x48));
  assign z27 = x53 & ~x52 & ~x51 & ~x50 & ~x49 & x48 & ~x46 & ~x47;
  assign z28 = ~x46 & x47 & ((x51 & ((x52 & ((~x48 & x50 & (x53 | (x49 & ~x53))) | (x49 & ~x50 & (~x53 | (x48 & x53))))) | (~x48 & x49 & ~x50 & ~x52 & x53))) | (~x48 & x49 & ~x50 & ~x51 & ~x52 & ~x53));
  assign z29 = x53 & ~x52 & x51 & x50 & x49 & x48 & ~x46 & x47;
  assign z30 = ~x47 & ((~x48 & ((~x51 & ((x49 & (x46 ? ((x52 & x53) | (x50 & ~x52 & ~x53)) : (~x50 & ~x52))) | (~x46 & ~x49 & x50 & (~x53 | (~x52 & x53))))) | (x46 & x49 & ~x50 & x51 & (x52 | (~x52 & (x24 | ~x53 | (~x24 & x53))))))) | (x46 & x48 & ~x49 & ~x50 & x51 & x52 & ~x53));
  assign z31 = ~x53 & x52 & x51 & ~x50 & x49 & ~x48 & ~x46 & ~x47;
  assign z32 = ~x47 & x49 & ((x51 & x52 & x53 & x46 & ~x48 & x50) | (~x51 & ~x52 & ~x53 & ~x46 & x48 & ~x50));
  assign z33 = ~x53 & ~x52 & x51 & x50 & x49 & x48 & ~x46 & x47;
  assign z34 = ~x46 & x47 & x49 & ~x50 & ~x51 & ((~x52 & (x53 | (x48 & ~x53))) | (~x48 & x52 & ~x53));
  assign z35 = (x49 & ((~x46 & x50 & ~x51 & x53 & (x47 ? (~x48 & ~x52) : (x48 & x52))) | (~x50 & x51 & x52 & ~x53 & x46 & ~x47 & ~x48))) | (~x46 & ~x47 & x48 & ~x49 & ~x53 & ((~x51 & x52) | (x50 & x51 & ~x52)));
  assign z36 = x53 & x52 & ~x51 & ~x50 & x49 & x48 & ~x46 & ~x47;
  assign z37 = ~x53 & ~x52 & ~x51 & ~x50 & x49 & x48 & ~x46 & ~x47;
  assign z38 = ~x53 & ~x52 & x51 & ~x50 & x49 & x48 & ~x46 & ~x47;
  assign z39 = ~x46 & ~x47 & x48 & ~x49 & ~x52 & x53 & ((~x50 & x51) | (~x24 & x50 & ~x51));
  assign z40 = ~x52 & ((~x51 & ((~x46 & x47 & x49 & x50 & (x48 | (~x48 & ~x53))) | (x46 & ~x47 & x48 & ~x49 & ~x50 & x53))) | (~x46 & x47 & ~x48 & x50 & (x53 ? x51 : (x49 ? (x11 | (~x11 & x51)) : x51))));
  assign z41 = ~x50 & ((x51 & x52 & x53 & ~x46 & x47 & ~x49) | (x46 & ~x47 & ~x48 & ~x52 & ~x53 & x49 & ~x51));
  assign z42 = x53 & x52 & x51 & ~x50 & x49 & ~x48 & ~x46 & ~x47;
  assign z43 = x53 & ~x52 & x51 & ~x50 & x49 & ~x48 & ~x46 & ~x47;
  assign z44 = ~x46 & ~x47 & x48 & ~x49 & ((x50 & (x51 ^ x52)) | (x52 & x53 & ~x50 & ~x51));
  assign z45 = ~x53 & x52 & x51 & ~x50 & x49 & ~x48 & ~x46 & ~x47;
  assign z46 = x53 & x52 & x51 & x50 & x49 & x48 & ~x46 & x47;
  assign z47 = ~x53 & ~x52 & x51 & ~x50 & ~x49 & x48 & ~x46 & ~x47;
  assign z48 = ~x53 & ~x52 & x51 & ~x50 & ~x49 & ~x48 & x47 & ~x46 & x27 & ~x43;
  assign z49 = (~x48 & ((~x50 & ((x51 & x52 & x53 & ~x46 & x47 & ~x49) | (~x47 & ((x46 & x49 & x52 & (x51 ^ x53)) | (x51 & ~x52 & x53 & ~x46 & ~x49))))) | (x52 & x53 & x50 & ~x51 & ~x46 & x47 & ~x49))) | (x52 & x53 & x50 & ~x51 & x46 & ~x47 & x48 & ~x49);
endmodule