module pla__shift ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15;
  assign z00 = x03;
  assign z01 = (x03 & ((x00 & (~x01 | (x01 & x02))) | (~x00 & x02) | (x01 & ~x02))) | (~x00 & ~x01 & ~x02 & x04);
  assign z02 = x01 ? x03 : (x00 ? x03 : (x02 ? x04 : x05));
  assign z03 = (x03 & ((x01 & x02) | (x00 & (~x01 | (x01 & ~x02))))) | (~x00 & (x01 ? (~x02 & x04) : (x02 ? x05 : x06)));
  assign z04 = x00 ? x03 : (x01 ? (x02 ? x04 : x05) : (x02 ? x06 : x07));
  assign z05 = x00 ? (x02 ? x03 : (x01 ? x03 : x04)) : (x01 ? (x02 ? x05 : x06) : (x02 ? x07 : x08));
  assign z06 = x01 ? (x00 ? x03 : (x02 ? x06 : x07)) : (x00 ? (x02 ? x04 : x05) : (x02 ? x08 : x09));
  assign z07 = x00 ? (x01 ? (x02 ? x03 : x04) : (x02 ? x05 : x06)) : (x01 ? (x02 ? x07 : x08) : (x02 ? x09 : x10));
  assign z08 = x00 ? (x01 ? (x02 ? x04 : x05) : (x02 ? x06 : x07)) : (x01 ? (x02 ? x08 : x09) : (x02 ? x10 : x11));
  assign z09 = x00 ? (x01 ? (x02 ? x05 : x06) : (x02 ? x07 : x08)) : (x01 ? (x02 ? x09 : x10) : (x02 ? x11 : x12));
  assign z10 = x00 ? (x01 ? (x02 ? x06 : x07) : (x02 ? x08 : x09)) : (x01 ? (x02 ? x10 : x11) : (x02 ? x12 : x13));
  assign z11 = x00 ? (x01 ? (x02 ? x07 : x08) : (x02 ? x09 : x10)) : (x01 ? (x02 ? x11 : x12) : (x02 ? x13 : x14));
  assign z12 = x00 ? (x01 ? (x02 ? x08 : x09) : (x02 ? x10 : x11)) : (x01 ? (x02 ? x12 : x13) : (x02 ? x14 : x15));
  assign z13 = x00 ? (x01 ? (x02 ? x09 : x10) : (x02 ? x11 : x12)) : (x01 ? (x02 ? x13 : x14) : (x02 ? x15 : x16));
  assign z14 = x00 ? (x01 ? (x02 ? x10 : x11) : (x02 ? x12 : x13)) : (x01 ? (x02 ? x14 : x15) : (x02 ? x16 : x17));
  assign z15 = x00 ? (x01 ? (x02 ? x11 : x12) : (x02 ? x13 : x14)) : (x01 ? (x02 ? x15 : x16) : (x02 ? x17 : x18));
endmodule