module pla__amd ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23;
  assign z00 = (x06 & ((~x10 & ((~x05 & ((~x00 & ((~x09 & x13) | (x04 & x09 & ~x11 & x12 & ~x13))) | (~x11 & ((x00 & ~x04 & (x09 ^ x13)) | (x04 & x09 & x12 & x13))) | (x00 & ~x09 & x11 & ~x12 & (~x13 | (~x04 & x13))))) | (~x03 & x05 & (x09 ? ~x11 : (x12 | (x11 & ~x12)))))) | (~x09 & ((~x11 & ((~x03 & x05 & (x13 ? ~x12 : x10)) | (x10 & ((x12 & x13) | (~x05 & (x00 ? (x12 & ~x13) : (~x12 & x13))))))) | (x10 & x11 & x13 & (~x12 | (x12 & (x01 | (~x01 & ~x03))))))))) | (~x05 & ((~x06 & ((x09 & ~x10 & ~x11 & x13) | (x08 & ~x09 & x10 & x11 & ~x12 & ~x13))) | (~x10 & ~x12 & ~x13 & ((x09 & x11) | (x03 & x08 & ~x09 & ~x11)))));
  assign z01 = (x06 & (x09 ? (~x10 & ~x11 & (x05 | (~x05 & ~x13 & (x00 ? (~x12 | (x04 & x12)) : x12)))) : ((~x05 & (x00 ? ((x10 & ~x11 & ~x13) | (x04 & ~x10 & x13 & (~x11 | (x11 & ~x12)))) : (x12 & (~x10 | (x10 & ~x11 & ~x13))))) | (x05 & ((~x10 & (x12 | (x11 & ~x12))) | (~x11 & (x13 ? ~x12 : x10)))) | (x10 & x12 & (x11 ? ~x01 : x13))))) | (~x05 & x09 & ~x10 & (x11 ? (~x12 & ~x13) : (x12 & x13)));
  assign z02 = (x06 & ((~x10 & (x05 ? (x09 ? ~x11 : (x12 | (x11 & ~x12))) : ((~x00 & ((x04 & x09 & ~x11 & x12 & ~x13) | (~x09 & x11))) | (~x11 & ((x00 & x12 & ~x13) | (x13 & ((x00 & ~x09 & (x04 | (~x04 & ~x12))) | (x04 & x09 & x12))))) | (x00 & ~x09 & x11 & (x12 | (~x12 & x13)))))) | (~x09 & ((x05 & ~x11 & (x13 ? ~x12 : x10)) | (x10 & x11))))) | (~x04 & ~x05 & ~x08 & ~x09 & ~x12 & ~x13 & ((~x06 & x10 & x11) | (x03 & ~x10 & ~x11)));
  assign z03 = x06 & ((~x09 & ((~x11 & ((x05 & (x13 ? ~x12 : x10)) | (x10 & ((x12 & x13) | (~x05 & (~x12 | (x12 & ~x13))))))) | (x10 & x11) | (~x10 & ((x05 & (x12 | (x11 & ~x12))) | (x11 & ~x12 & ~x13 & x00 & ~x05))))) | (~x10 & ~x11 & x05 & x09));
  assign z04 = ~x05 & ((~x10 & ((~x11 & ((x09 & (x06 ? ((~x12 | (~x04 & x12)) & (x13 | (~x00 & ~x13))) : x13)) | (x03 & ~x09 & ~x12 & ~x13 & (~x04 | (x04 & x08))))) | (~x12 & ~x13 & x09 & x11))) | (~x06 & ~x09 & x10 & x11 & ~x12 & ~x13 & (~x04 | (x04 & x08))));
  assign z05 = ~x05 & ~x09 & ~x12 & ~x13 & ((~x06 & x10 & x11) | (x03 & ~x10 & ~x11));
  assign z06 = x00 & x02 & ~x05 & x06 & ~x10 & ((~x09 & (x12 ? x11 : x13)) | (x12 & ~x13 & x09 & ~x11));
  assign z07 = x07 & ((~x09 & (x06 ? ((~x05 & ((~x11 & (x00 ? (x12 ? ~x13 : x10) : (x13 ? ~x12 : x10))) | (~x10 & (x00 ? (x13 | (x11 & ~x13)) : (x12 | (x11 & ~x12)))))) | (x10 & ((x11 & x12) | (x05 & ~x11 & ~x13))) | (x05 & ((~x10 & (x12 | (x11 & ~x12))) | (~x11 & ~x12 & x13)))) : ((~x10 & (~x11 ^ ~x12)) | (~x11 & (x13 ? ~x12 : x10)) | (x11 & x12)))) | (x09 & ~x10 & ~x11 & ~x13));
  assign z08 = x13 & ~x12 & x11 & x10 & ~x06 & ~x09;
  assign z09 = x13 & x12 & ~x11 & x10 & ~x06 & ~x09;
  assign z10 = ~x05 & ~x10 & ((x09 & ~x13 & ((x11 & ~x12) | (~x11 & x12 & x00 & x06))) | (x00 & x06 & ~x09 & x13 & (~x11 | (x11 & ~x12))));
  assign z11 = x00 & ~x05 & x06 & ~x10 & ((x12 & x13 & ~x09 & x11) | (x09 & ~x11 & ~x13));
  assign z12 = x05 ? (x06 & (x09 ? (~x10 & ~x11) : ((~x10 & (x12 | (x11 & ~x12))) | (~x11 & (x13 ? ~x12 : x10))))) : ((~x06 & ((x09 & ~x10 & ~x11 & x13) | (x08 & ~x09 & x10 & x11 & ~x12 & ~x13))) | (~x10 & ~x12 & ~x13 & ((x09 & x11) | (x03 & x08 & ~x09 & ~x11))));
  assign z13 = x05 & x06 & (x09 ? (~x10 & ~x11) : ((~x10 & (x12 | (x11 & ~x12))) | (~x11 & (x13 ? ~x12 : x10))));
  assign z14 = ~x05 & ((~x06 & ((x09 & ~x10 & ~x11 & x13) | (x08 & ~x09 & x10 & x11 & ~x12 & ~x13))) | (~x12 & ~x13 & (x09 ? (~x10 & x11) : (~x11 & ((x00 & x06 & x10) | (x03 & x08 & ~x10))))));
  assign z15 = x12 & ~x11 & ~x10 & ~x09 & x06 & x00 & ~x05;
  assign z16 = ~x13 & ~x12 & ~x11 & ~x10 & x09 & x06 & x00 & ~x05;
  assign z17 = x00 & ~x05 & x06 & ~x10 & ((~x09 & (x12 ? x11 : x13)) | (x12 & ~x13 & x09 & ~x11));
  assign z18 = x05 ? (x06 & (x09 ? (~x10 & ~x11) : ((~x10 & (x12 | (x11 & ~x12))) | (~x11 & (x13 ? ~x12 : x10))))) : ((~x06 & ((x09 & ~x10 & ~x11 & x13) | (x08 & ~x09 & x10 & x11 & ~x12 & ~x13))) | (~x10 & ((~x13 & ((x09 & ((x11 & ~x12) | (x00 & x06 & ~x11))) | (x03 & x08 & ~x09 & ~x11 & ~x12))) | (x00 & x06 & ~x09 & (x12 | (~x12 & x13))))) | (x00 & x06 & ~x09 & ~x12 & ~x13 & x10 & ~x11));
  assign z19 = ~x05 & ((~x10 & ((x06 & ((~x09 & x13 & (~x11 | (x11 & ~x12)) & (~x00 | (x00 & ~x04))) | (~x04 & x09 & ~x11 & (x12 | (x00 & ~x12 & ~x13))))) | (x09 & ((x11 & ~x12 & ~x13) | (x12 & x13 & ~x06 & ~x11))) | (x03 & ~x04 & ~x08 & ~x12 & ~x13 & ~x09 & ~x11))) | (~x04 & ~x06 & ~x08 & ~x09 & ~x12 & ~x13 & x10 & x11));
  assign z20 = ~x04 & ~x05 & ~x08 & ~x09 & ~x12 & ~x13 & ((~x06 & x10 & x11) | (x03 & ~x10 & ~x11));
  assign z21 = ~x05 & x06 & ((~x09 & ((~x10 & (x12 ? ((x00 & (x13 | (~x11 & ~x13))) | (x11 & ~x13) | (~x00 & ~x11)) : x11)) | (~x11 & ~x12 & (x13 | (~x00 & x10 & ~x13))))) | (x00 & x09 & ~x10 & ~x11 & ~x13));
  assign z22 = ~x05 & x06 & ~x09 & ~x12 & ((x10 & ~x11 & (x13 | (~x00 & ~x13))) | (x11 & ~x13 & x00 & ~x10));
  assign z23 = (x06 & (x09 ? (~x10 & ~x11 & (x05 | (~x05 & ~x13))) : ((~x11 & (x05 ? (x13 ? ~x12 : x10) : ((~x00 & x10 & ~x13) | (~x12 & (x00 ? (x10 | (~x10 & x13)) : x13))))) | (~x10 & (x12 | (x11 & ~x12))) | (x11 & x12 & ~x01 & x10)))) | (~x05 & ((x09 & ~x10 & ~x11 & x13) | (~x12 & ~x13 & ((x09 & ~x10 & x11) | (x08 & ~x09 & ((~x06 & x10 & x11) | (x03 & ~x10 & ~x11)))))));
endmodule