module pla__o64 ( 
    x000, x001, x002, x003, x004, x005, x006, x007, x008, x009, x010, x011,
    x012, x013, x014, x015, x016, x017, x018, x019, x020, x021, x022, x023,
    x024, x025, x026, x027, x028, x029, x030, x031, x032, x033, x034, x035,
    x036, x037, x038, x039, x040, x041, x042, x043, x044, x045, x046, x047,
    x048, x049, x050, x051, x052, x053, x054, x055, x056, x057, x058, x059,
    x060, x061, x062, x063, x064, x065, x066, x067, x068, x069, x070, x071,
    x072, x073, x074, x075, x076, x077, x078, x079, x080, x081, x082, x083,
    x084, x085, x086, x087, x088, x089, x090, x091, x092, x093, x094, x095,
    x096, x097, x098, x099, x100, x101, x102, x103, x104, x105, x106, x107,
    x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119,
    x120, x121, x122, x123, x124, x125, x126, x127, x128, x129,
    z0  );
  input  x000, x001, x002, x003, x004, x005, x006, x007, x008, x009,
    x010, x011, x012, x013, x014, x015, x016, x017, x018, x019, x020, x021,
    x022, x023, x024, x025, x026, x027, x028, x029, x030, x031, x032, x033,
    x034, x035, x036, x037, x038, x039, x040, x041, x042, x043, x044, x045,
    x046, x047, x048, x049, x050, x051, x052, x053, x054, x055, x056, x057,
    x058, x059, x060, x061, x062, x063, x064, x065, x066, x067, x068, x069,
    x070, x071, x072, x073, x074, x075, x076, x077, x078, x079, x080, x081,
    x082, x083, x084, x085, x086, x087, x088, x089, x090, x091, x092, x093,
    x094, x095, x096, x097, x098, x099, x100, x101, x102, x103, x104, x105,
    x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117,
    x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129;
  output z0;
  assign z0 = (x000 & x129) | (x064 & x128) | (x063 & x127) | (x062 & x126) | (x061 & x125) | (x060 & x124) | (x059 & x123) | (x058 & x122) | (x057 & x121) | (x056 & x120) | (x055 & x119) | (x054 & x118) | (x053 & x117) | (x052 & x116) | (x051 & x115) | (x050 & x114) | (x049 & x113) | (x048 & x112) | (x047 & x111) | (x046 & x110) | (x045 & x109) | (x044 & x108) | (x043 & x107) | (x042 & x106) | (x041 & x105) | (x040 & x104) | (x039 & x103) | (x038 & x102) | (x037 & x101) | (x036 & x100) | (x035 & x099) | (x034 & x098) | (x033 & x097) | (x032 & x096) | (x031 & x095) | (x030 & x094) | (x029 & x093) | (x028 & x092) | (x027 & x091) | (x026 & x090) | (x025 & x089) | (x024 & x088) | (x023 & x087) | (x022 & x086) | (x021 & x085) | (x020 & x084) | (x019 & x083) | (x018 & x082) | (x017 & x081) | (x016 & x080) | (x015 & x079) | (x014 & x078) | (x013 & x077) | (x012 & x076) | (x011 & x075) | (x010 & x074) | (x009 & x073) | (x008 & x072) | (x007 & x071) | (x006 & x070) | (x005 & x069) | (x004 & x068) | (x003 & x067) | (x002 & x066) | (x001 & x065);
endmodule