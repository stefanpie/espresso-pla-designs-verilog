module pla__dk17 ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10;
  assign z00 = ~x1 & ~x3 & ~x4 & ~x5 & ~x7 & ~x8 & ((~x0 & (x2 ? ~x6 : (x6 & x9))) | (x0 & ~x2 & ~x6 & ~x9));
  assign z01 = ~x1 & ~x3 & ~x4 & ~x5 & ~x7 & x8 & ((~x0 & (x2 ? ~x6 : (x6 & x9))) | (x0 & ~x2 & ~x6 & ~x9));
  assign z02 = ~x0 & ~x2 & ~x3 & ~x6 & ((~x1 & ((~x5 & (x4 ? (~x7 & (~x9 | (x8 & x9))) : (x7 & x8))) | (~x4 & x5 & ~x7 & x8))) | (x1 & ~x4 & ~x5 & ~x7 & ~x9));
  assign z03 = ~x2 & ~x5 & ((~x0 & ((~x3 & ~x8 & ((~x6 & ((~x1 & (x4 ? (~x7 & x9) : (x7 & ~x9))) | (x1 & ~x4 & ~x7 & x9))) | (~x1 & ~x4 & x6 & ~x7 & ~x9))) | (~x1 & x3 & ~x4 & ~x6 & ~x7 & ~x9))) | (x0 & ~x1 & ~x3 & ~x4 & ~x6 & ~x7 & ~x8 & x9));
  assign z04 = ~x1 & ~x2 & ~x4 & ~x5 & ((~x3 & ((~x0 & ((~x8 & x9 & ~x6 & x7) | (x6 & ~x7 & x8 & ~x9))) | (x0 & ~x6 & ~x7 & x8 & x9))) | (~x0 & x3 & ~x6 & ~x7 & x9));
  assign z05 = x9 & x8 & ~x7 & ~x6 & ~x5 & ~x4 & ~x3 & ~x2 & ~x0 & x1;
  assign z06 = ~x9 & ~x8 & ~x7 & ~x6 & x5 & ~x4 & ~x3 & ~x2 & ~x0 & ~x1;
  assign z07 = x9 & ~x8 & ~x7 & ~x6 & x5 & ~x4 & ~x3 & ~x2 & ~x0 & ~x1;
  assign z08 = ~x0 & ~x1 & ((~x2 & ((~x3 & ((~x4 & ((~x5 & (x6 ? (~x7 & x9) : (x7 & (~x8 | (x8 & x9))))) | (~x7 & x8 & x9 & x5 & ~x6))) | (~x7 & x8 & x9 & x4 & ~x5 & ~x6))) | (x3 & ~x4 & ~x5 & ~x6 & ~x7 & ~x8))) | (x2 & ~x3 & ~x4 & ~x7 & x9 & ~x5 & ~x6));
  assign z09 = ~x2 & ((~x0 & ((~x1 & ((~x3 & ~x9 & ((~x4 & ((~x5 & (x6 ? ~x7 : (x7 & x8))) | (~x7 & x8 & x5 & ~x6))) | (x4 & ~x5 & ~x6 & ~x7 & x8))) | (x3 & ~x4 & ~x5 & ~x6 & ~x7 & x8))) | (~x4 & ~x5 & x1 & ~x3 & ~x6 & ~x7 & x8 & ~x9))) | (x0 & ~x1 & ~x3 & ~x4 & ~x7 & x9 & ~x5 & ~x6));
  assign z10 = ~x1 & ~x3 & ~x4 & ~x5 & ~x7 & ((~x0 & (x2 ? ~x6 : (x6 & x9))) | (x0 & ~x2 & ~x6 & ~x9));
endmodule