module pla__newcpla2 ( 
    CPIPE2s__larrow__0__rarrow__, CPIPE2s__larrow__1__rarrow__,
    CPIPE2s__larrow__2__rarrow__, CPIPE2s__larrow__3__rarrow__,
    CPIPE2s__larrow__4__rarrow__, CPIPE2s__larrow__5__rarrow__,
    CPIPE2s__larrow__7__rarrow__,
    writeRFaccess2, lastPCtobusD1, busDtobusB2, busDtobusA2, DSTtobusD2,
    nillonreturn, pLOADwrite, opc2load, DSTvalid, pbusDtoINA  );
  input  CPIPE2s__larrow__0__rarrow__, CPIPE2s__larrow__1__rarrow__,
    CPIPE2s__larrow__2__rarrow__, CPIPE2s__larrow__3__rarrow__,
    CPIPE2s__larrow__4__rarrow__, CPIPE2s__larrow__5__rarrow__,
    CPIPE2s__larrow__7__rarrow__;
  output writeRFaccess2, lastPCtobusD1, busDtobusB2, busDtobusA2, DSTtobusD2,
    nillonreturn, pLOADwrite, opc2load, DSTvalid, pbusDtoINA;
  assign writeRFaccess2 = (CPIPE2s__larrow__7__rarrow__ & ((~CPIPE2s__larrow__2__rarrow__ & ((~CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__4__rarrow__) | (CPIPE2s__larrow__0__rarrow__ & CPIPE2s__larrow__3__rarrow__ & CPIPE2s__larrow__4__rarrow__ & ~CPIPE2s__larrow__5__rarrow__))) | (CPIPE2s__larrow__1__rarrow__ & ((CPIPE2s__larrow__0__rarrow__ & (~CPIPE2s__larrow__4__rarrow__ | (CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__))) | (CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__4__rarrow__ & ~CPIPE2s__larrow__5__rarrow__))) | (CPIPE2s__larrow__5__rarrow__ & (~CPIPE2s__larrow__4__rarrow__ | (~CPIPE2s__larrow__3__rarrow__ & CPIPE2s__larrow__4__rarrow__))))) | (~CPIPE2s__larrow__5__rarrow__ & (~CPIPE2s__larrow__7__rarrow__ | (CPIPE2s__larrow__0__rarrow__ & ~CPIPE2s__larrow__1__rarrow__ & CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__4__rarrow__)));
  assign lastPCtobusD1 = ~CPIPE2s__larrow__5__rarrow__ & (~CPIPE2s__larrow__7__rarrow__ | (CPIPE2s__larrow__0__rarrow__ & ~CPIPE2s__larrow__1__rarrow__ & CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__4__rarrow__));
  assign busDtobusB2 = (~CPIPE2s__larrow__4__rarrow__ & ((CPIPE2s__larrow__7__rarrow__ & ((CPIPE2s__larrow__1__rarrow__ & ((CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__) | (CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & CPIPE2s__larrow__5__rarrow__))) | (CPIPE2s__larrow__5__rarrow__ & (~CPIPE2s__larrow__0__rarrow__ | (~CPIPE2s__larrow__1__rarrow__ & ~CPIPE2s__larrow__2__rarrow__ & CPIPE2s__larrow__3__rarrow__))))) | (CPIPE2s__larrow__0__rarrow__ & ~CPIPE2s__larrow__1__rarrow__ & CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__))) | (~CPIPE2s__larrow__5__rarrow__ & ~CPIPE2s__larrow__7__rarrow__);
  assign busDtobusA2 = (~CPIPE2s__larrow__4__rarrow__ & ((CPIPE2s__larrow__7__rarrow__ & ((CPIPE2s__larrow__1__rarrow__ & ((CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__) | (CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & CPIPE2s__larrow__5__rarrow__))) | (CPIPE2s__larrow__5__rarrow__ & (~CPIPE2s__larrow__0__rarrow__ | (~CPIPE2s__larrow__1__rarrow__ & ~CPIPE2s__larrow__2__rarrow__ & CPIPE2s__larrow__3__rarrow__))))) | (CPIPE2s__larrow__0__rarrow__ & ~CPIPE2s__larrow__1__rarrow__ & CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__))) | (~CPIPE2s__larrow__5__rarrow__ & ~CPIPE2s__larrow__7__rarrow__);
  assign DSTtobusD2 = ~CPIPE2s__larrow__4__rarrow__ & CPIPE2s__larrow__7__rarrow__ & ((CPIPE2s__larrow__1__rarrow__ & ((CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__) | (CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & CPIPE2s__larrow__5__rarrow__))) | (CPIPE2s__larrow__5__rarrow__ & (~CPIPE2s__larrow__0__rarrow__ | (~CPIPE2s__larrow__1__rarrow__ & ~CPIPE2s__larrow__2__rarrow__ & CPIPE2s__larrow__3__rarrow__))));
  assign nillonreturn = CPIPE2s__larrow__7__rarrow__ & ~CPIPE2s__larrow__5__rarrow__ & ~CPIPE2s__larrow__4__rarrow__ & CPIPE2s__larrow__1__rarrow__ & CPIPE2s__larrow__3__rarrow__;
  assign pLOADwrite = CPIPE2s__larrow__7__rarrow__ & CPIPE2s__larrow__5__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & CPIPE2s__larrow__4__rarrow__;
  assign opc2load = CPIPE2s__larrow__7__rarrow__ & CPIPE2s__larrow__5__rarrow__ & CPIPE2s__larrow__4__rarrow__ & ~CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__2__rarrow__ & ~CPIPE2s__larrow__0__rarrow__ & ~CPIPE2s__larrow__1__rarrow__;
  assign DSTvalid = CPIPE2s__larrow__7__rarrow__ & ((CPIPE2s__larrow__0__rarrow__ & ((CPIPE2s__larrow__1__rarrow__ & (~CPIPE2s__larrow__4__rarrow__ | (CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__))) | (CPIPE2s__larrow__4__rarrow__ & ~CPIPE2s__larrow__5__rarrow__ & ~CPIPE2s__larrow__2__rarrow__ & CPIPE2s__larrow__3__rarrow__))) | (~CPIPE2s__larrow__3__rarrow__ & (CPIPE2s__larrow__4__rarrow__ ? CPIPE2s__larrow__5__rarrow__ : ~CPIPE2s__larrow__2__rarrow__)) | (~CPIPE2s__larrow__4__rarrow__ & (CPIPE2s__larrow__3__rarrow__ | CPIPE2s__larrow__5__rarrow__)));
  assign pbusDtoINA = CPIPE2s__larrow__4__rarrow__ & CPIPE2s__larrow__7__rarrow__ & ((CPIPE2s__larrow__2__rarrow__ & (CPIPE2s__larrow__5__rarrow__ | (~CPIPE2s__larrow__1__rarrow__ & CPIPE2s__larrow__3__rarrow__))) | (CPIPE2s__larrow__5__rarrow__ & (CPIPE2s__larrow__0__rarrow__ | CPIPE2s__larrow__1__rarrow__)) | (~CPIPE2s__larrow__0__rarrow__ & CPIPE2s__larrow__3__rarrow__ & ~CPIPE2s__larrow__5__rarrow__));
endmodule