module pla__in3 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28;
  assign z00 = x00 ? ((~x03 & (x01 ? (~x02 & ((~x17 & ((~x06 & ~x07 & x08 & (x25 | (~x09 & ~x25 & ~x33 & ~x34))) | (~x34 & (x33 | (x06 & ~x33))))) | (x17 & (~x28 | (x28 & (~x26 | (x26 & ~x34))))) | x34 | (~x33 & ~x34 & x08 & x09))) : (x02 & (~x29 | (x29 & x30))))) | (~x01 & x02 & (~x30 | (x03 & x30)))) : ((x01 & x02 & x03) | (~x01 & ~x02 & ~x03 & x22 & ~x34));
  assign z01 = (x02 & ((~x01 & (~x00 | (x00 & x03 & x30))) | (~x00 & x01 & (x03 ? (x08 | (~x08 & x17)) : (~x34 & (x17 | (~x17 & ~x33 & ((~x06 & (x09 | (~x09 & (x10 | (~x07 & ~x08 & (x27 | (~x27 & ~x32))))))) | x06 | (~x07 & x08))))))))) | (x01 & ~x02 & (~x00 | (x00 & ~x03 & ((x17 & (~x28 | (~x26 & x28))) | x34 | (~x17 & ((~x06 & ~x07 & x08 & x25) | (x33 & ~x34)))))));
  assign z02 = (~x03 & ((~x34 & ((x01 & ((~x33 & ((~x17 & (x00 ? (~x02 & (x06 | (~x06 & ~x07 & x08 & ~x09 & ~x25))) : (x02 & ((~x06 & (x09 | (~x09 & (x10 | (~x07 & ~x08 & (x27 | (~x27 & ~x32))))))) | x06 | (~x07 & x08))))) | (x08 & x09 & x00 & ~x02))) | (x17 & ((~x00 & x02) | (x00 & ~x02 & x26 & x28))))) | (~x00 & ~x01 & ~x02 & x22))) | (~x01 & (x00 ? (x02 & (~x29 | (x29 & x30))) : (~x02 & ~x22 & x29 & (x21 | (x20 & ~x21))))))) | (x00 & ~x01 & x02 & (~x30 | (x03 & x30))) | (~x00 & x01 & ~x02 & x30);
  assign z03 = x01 ? (~x03 & ((~x17 & (x00 ? (~x02 & ((~x06 & ~x07 & x08 & x25) | (x33 & ~x34))) : (x02 & ~x33 & ~x34 & ((~x06 & (x09 | (~x09 & (x10 | (~x07 & ~x08 & (x27 | (~x27 & ~x32))))))) | x06 | (~x07 & x08))))) | (x00 & ~x02 & (x34 | (x17 & (~x28 | (~x26 & x28))))) | (~x00 & x02 & x17 & ~x34))) : ((x00 & (x02 ? (x03 ? ~x30 : (x29 & x30)) : ~x03)) | (~x02 & x03 & x10));
  assign z04 = ~x00 & x01 & x02 & ~x03 & ~x17 & ~x18 & x24 & ~x27 & x32 & ~x33 & ~x34 & (~x14 | (x04 & ~x05 & x14));
  assign z05 = (x01 & (x00 ? (x02 ? ~x19 : x03) : ((x02 & ~x03 & (x34 | (~x17 & ~x34 & (x33 | (x24 & ~x27 & x32 & ~x33 & (x18 | (x14 & ~x18 & (~x04 | (x04 & x05))))))))) | (~x02 & ~x06 & ~x07 & ~x08 & x30)))) | (~x01 & ~x02 & x03 & ~x10);
  assign z06 = x19 & x02 & x00 & x01;
  assign z07 = ~x00 & ~x01 & (x02 | (x22 & ~x34 & ~x02 & ~x03));
  assign z08 = (~x01 & ((x00 & x02) | (~x03 & x22 & ~x34 & ~x00 & ~x02))) | (x00 & x01 & ~x02 & ~x03 & ~x34 & ((~x33 & ((x08 & (x09 | (~x06 & ~x07 & ~x09 & ~x17 & ~x25))) | (x06 & ~x17))) | (x17 & x26 & x28)));
  assign z09 = (~x00 & x01 & ~x02 & x30) | (x00 & ~x01 & x02 & (x03 | (~x03 & x29 & x30)));
  assign z10 = (x00 & x01 & ~x02 & ~x03 & ~x34 & ((~x33 & ((x08 & (x09 | (~x06 & ~x07 & ~x09 & ~x17 & ~x25))) | (x06 & ~x17))) | (x17 & x26 & x28))) | (~x01 & ((~x03 & x22 & ~x34 & ~x00 & ~x02) | (x02 & (~x00 | (x00 & ~x03 & (~x29 | ~x30))))));
  assign z11 = ~x00 & ~x01 & ~x02 & ~x03 & ~x22 & x29 & (x21 | (x20 & ~x21));
  assign z12 = x00 ? ((~x03 & (x01 ? (~x02 & ~x34 & ((~x33 & ((x08 & (x09 | (~x06 & ~x07 & ~x09 & ~x17 & ~x25))) | (x06 & ~x17))) | (x17 & x26 & x28))) : (x02 & (~x29 | (x29 & x30 & ~x31))))) | (~x01 & x02 & ~x30)) : (x01 ? (((x08 | (~x08 & x17)) & (~x02 | (x02 & x03))) | (x02 & ~x03 & ~x34 & (x17 | (~x17 & ~x33 & (x08 | (~x18 & x24 & ~x27 & x32 & (~x14 | (x04 & ~x05 & x14)))))))) : (x02 ? (x17 | (x08 & ~x17)) : (~x03 & (x22 ? ~x34 : (x21 | (x20 & ~x21))))));
  assign z13 = ~x02 & ~x03 & ~x34 & (x00 ? (x01 & ((~x33 & ((x08 & (x09 | (~x06 & ~x07 & ~x09 & ~x17 & ~x25))) | (x06 & ~x17))) | (x17 & x26 & x28))) : (~x01 & x22));
  assign z14 = x01 ? ((x03 & ((x00 & ~x02) | (~x00 & x02 & ~x08 & ~x17))) | (~x03 & (x00 ? (~x02 & ((x17 & (~x28 | (~x26 & x28))) | x34 | (~x17 & ((~x06 & ~x07 & x08 & x25) | (x33 & ~x34))))) : (x02 & (x34 | (~x34 & ((~x17 & (x33 | (x24 & ~x27 & x32 & ~x33))) | (~x08 & ~x33))))))) | (x00 & x02) | (~x00 & ~x02)) : (~x02 | (~x00 & x02));
  assign z15 = (x03 & ((~x00 & x01 & x02) | (~x01 & ~x02 & x10))) | (x01 & ((~x03 & ~x34 & ((x17 & ((~x00 & x02) | (x00 & ~x02 & x26 & x28))) | (~x33 & ((x08 & x09 & x00 & ~x02) | (~x17 & (x00 ? (~x02 & (x06 | (~x06 & ~x07 & x08 & ~x09 & ~x25))) : (x02 & ((~x06 & (x09 | (~x09 & (x10 | (~x07 & ~x08 & (x27 | (~x27 & ~x32))))))) | x06 | (~x07 & x08) | (~x18 & x24 & ~x27 & x32 & (~x14 | (x04 & ~x05 & x14))))))))))) | (~x00 & ~x02 & (x08 | ~x30 | (x30 & (x27 | ~x32 | (x07 & ~x27))))))) | (~x01 & (x02 | (~x02 & ~x03 & (x00 | (~x00 & ~x22 & (x21 | (x20 & ~x21)))))));
  assign z16 = x00 & x06 & ~x17 & ((~x01 & x02) | (x01 & ~x02 & ~x03 & ~x33 & ~x34));
  assign z17 = ~x00 & x01 & x02 & x03 & (x08 | (~x08 & (x17 | (~x09 & ~x17))));
  assign z18 = ~x00 & x01 & x02 & ~x03 & (x34 | (~x34 & (x17 ? x28 : (x33 | (~x33 & ((~x06 & (x09 | (~x07 & ~x08 & ~x09 & (x27 | (~x27 & ~x32))))) | x06 | (~x07 & x08) | (x24 & ~x27 & x32)))))));
  assign z19 = (~x01 & ~x02 & x03 & ~x10) | (x01 & (x00 ? (x02 | (~x02 & x03)) : (x02 & ~x03 & (x34 | (~x17 & ~x34 & (x33 | (x24 & ~x27 & x32 & ~x33 & (x18 | (x14 & ~x18 & (~x04 | (x04 & x05)))))))))));
  assign z20 = ~x00 & ~x03 & ((x01 & x02 & ~x17 & ~x18 & x24 & ~x27 & x32 & ~x33 & ~x34 & (~x14 | (x04 & ~x05 & x14))) | (~x01 & ~x02 & x21 & ~x22 & ~x29));
  assign z21 = x30 & ~x08 & ~x07 & ~x06 & ~x02 & ~x00 & x01;
  assign z22 = x01 ? (~x02 & ((~x17 & ((x00 & ~x03 & ((~x06 & ~x07 & x08 & x25) | (x33 & ~x34))) | (~x00 & ~x06 & ~x07 & ~x08 & x16 & ~x27 & x29 & ~x30 & x32))) | (x00 & ~x03 & x34))) : ((~x17 & x30 & ((x02 & ((x00 & ~x03 & x14 & ~x19 & x29) | (~x00 & ~x06 & ~x07 & ~x08 & ~x27 & x32 & x16 & ~x23))) | (~x00 & ~x02 & ~x03 & ~x06 & ~x07 & ~x08 & ~x14 & x16 & ~x22 & ~x27 & x29 & x32 & ((~x12 & ((~x11 & (x20 | (~x20 & x21))) | (~x20 & x21 & x11 & ~x15))) | (~x15 & x20))))) | (~x02 & ((x00 & ~x03 & (x10 | (~x07 & ~x10 & x16))) | (x03 & x07 & x16))));
  assign z23 = x34 & ~x21 & ~x20 & ~x03 & ~x02 & ~x00 & ~x01;
  assign z24 = (x00 & ~x01 & x02 & (~x30 | (~x03 & ~x29))) | (~x00 & x01 & ~x02 & x29 & ~x30);
  assign z25 = (~x01 & ~x03 & (x00 ? (x02 & (~x29 | ~x30)) : (~x02 & ~x22 & ~x29 & (x21 | (x20 & ~x21))))) | (~x00 & x01 & ~x02 & ~x29 & ~x30);
  assign z26 = ~x34 & ~x33 & x32 & ~x27 & x24 & ~x18 & ~x17 & x14 & ~x05 & x04 & ~x03 & x02 & ~x00 & x01;
  assign z27 = x00 & x01 & (x02 ? (x17 & ~x19) : x03);
  assign z28 = (~x01 & ~x02 & x03 & ~x10) | (x01 & (x00 ? (x02 | (~x02 & x03)) : ((x02 & ~x03 & (x34 | (~x17 & ~x34 & (x33 | (x24 & ~x27 & x32 & ~x33 & (x18 | (~x18 & (~x14 | (x14 & (~x04 | (x04 & x05))))))))))) | (~x02 & ~x06 & ~x07 & ~x08 & ~x27 & x32))));
endmodule