module pla__chkn ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28,
    z0, z1, z2, z3, z4, z5, z6  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28;
  output z0, z1, z2, z3, z4, z5, z6;
  assign z0 = ~x04 & x12 & x15 & ((x02 & x11 & x13 & x14 & x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & x23 & (~x24 | ~x26)) | (~x11 & (~x13 | ~x16)));
  assign z1 = ~x04 & x16 & ((~x11 & ~x15 & (x12 | ~x14)) | (~x02 & x11 & x12 & x13 & x14 & x15 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & ~x22 & x23 & x26));
  assign z2 = x03 & ~x04 & ((x14 & ((x11 & ((x13 & x16 & (x12 ? (x15 & ~x17 & ~x18 & ~x19 & ~x20 & x21 & x22 & ~x23 & ~x24 & ((~x02 & (~x25 | ~x26)) | (~x25 & ~x26))) : (x02 | ~x15))) | (~x12 & ~x13 & x15))) | (x02 & ~x11 & ~x12 & ~x13 & (~x15 | x16)))) | (~x11 & ~x14 & ((x02 & x13 & (x12 ? (x15 & x16) : ~x15)) | (~x12 & ~x15 & x16))));
  assign z3 = x10 & ((~x04 & ((x12 & ((x05 & (((~x09 | x11) & (~x13 | ~x15 | ~x16)) | (x11 & x14 & ~x17 & ~x18 & ~x19 & ~x20 & ((~x21 & ((~x02 & ((~x25 & ((x22 & (x23 | (~x24 & ~x26))) | (~x22 & ~x23 & ~x24 & x26))) | (~x09 & ~x22 & x23))) | (x23 & ((x02 & ((~x09 & (~x24 | ~x26)) | (x22 & ~x26))) | (x22 & ~x24))) | (~x23 & x24 & ((x02 & (x26 ? ~x22 : x25)) | (~x09 & x22 & (~x25 | x26)))))) | (~x22 & ((~x24 & ((x02 & (x21 | (~x09 & ~x25 & x26))) | (x21 & (x23 ? (x25 & x26) : ~x26)))) | (~x23 & x24 & x25 & (x02 | x21 | x26)))))))) | (x07 & ((~x15 & (x11 | ~x16)) | (x11 & ((x13 & x14 & ~x17 & ~x18 & ~x19 & ~x20 & ((~x22 & ((x23 & ((~x02 & ~x21 & ~x26) | (x25 & x26 & x21 & ~x24))) | (~x23 & ((x16 & (x02 ? ((x24 & x25) | (~x21 & ~x25 & x26)) : (~x21 & x25 & (~x24 | x26)))) | (~x26 & ((x21 & (x02 | ~x24)) | (~x24 & ~x25))) | (x21 & x24 & x25))) | (x02 & x21 & ~x24))) | (~x21 & ((~x02 & ((x22 & ((x23 & (~x24 | ~x25)) | (x25 & ~x26 & ~x23 & x24))) | (~x25 & ~x26 & ~x23 & ~x24))) | (x22 & x23 & ((~x24 & ~x25) | (x02 & ~x26))))))) | ~x16 | (~x13 & ~x14))))) | (x06 & x11 & x13 & x14 & x15 & x16 & ~x17 & ~x18 & ~x19 & ~x20 & ((~x22 & ((~x02 & ((~x21 & x25 & (~x24 | x26)) | (x23 & (~x21 | (~x24 & x25 & x26))))) | (~x23 & ((x02 & ~x21 & x26 & (x24 | ~x25)) | (x21 & ~x26 & (~x24 | x25)))) | (~x24 & ~x26 & x02 & x21))) | (~x21 & ((x23 & ((x02 & (~x24 | ~x26)) | (~x24 & ~x26) | (~x02 & ~x25))) | (x22 & ((~x23 & x24 & (~x25 | ~x26)) | (~x02 & ~x25 & ~x26))))))))) | (~x12 & ((~x14 & ((x05 & ~x09 & (x11 ? x13 : x16)) | (x07 & x15 & ((~x11 & (~x13 | x16)) | (~x13 & ~x16))) | (x08 & x11 & ~x13 & ~x15))) | (x13 & ((x05 & ((~x11 & (x14 | (x15 & x16))) | (x14 & x15 & ~x16))) | (~x11 & x14 & (x07 | (x06 & ~x16))))))) | (x05 & ~x09 & ~x11 & x15 & (x14 ? ~x16 : ~x13)) | (x07 & x13 & x14 & ~x15 & ~x16))) | (x07 & (x27 | x28)));
  assign z4 = x00 & ~x04 & ((x14 & x15 & ((~x09 & ((~x13 & ~x16 & ~x11 & ~x12) | (x11 & x12 & x13 & x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & x22 & ~x23 & x24))) | (x11 & x12 & x13 & x16 & ~x17 & ~x18 & ~x19 & ~x20 & ~x21 & x22 & ~x23 & ((x24 & (~x25 | ~x26)) | (~x02 & ~x25 & ~x26))))) | (x11 & ~x12 & (~x14 | ~x15 | (x13 & ~x16))));
  assign z5 = x01 & ~x04 & ((x14 & ((~x13 & ((~x11 & (~x15 | x16)) | (~x03 & x11 & ~x12 & x15))) | (x11 & x13 & x16 & ((~x12 & (~x03 | x15)) | (x15 & ~x17 & ~x18 & ~x19 & ~x20 & (((~x02 | ~x26) & ((~x22 & x23 & x24) | (~x03 & x21 & x22 & ~x23 & ~x24 & ~x25))) | (~x24 & ((~x21 & ~x22 & x23) | (~x02 & ~x03 & x21 & x22 & ~x23 & ~x26))))))))) | (~x11 & ((x12 & (~x14 | ~x15 | ~x16)) | (~x14 & ~x15 & (x13 | x16)))));
  assign z6 = ((~x13 | ~x15 | ~x16) & (x11 | x12)) | (~x12 & (x11 | x14 | x16)) | (x11 & x14 & ~x17 & ~x18 & ~x19 & ~x20 & ((~x21 & ((x22 & ((~x23 & x24) | (~x02 & ~x25 & ~x26))) | (x02 & (x23 ? ~x26 : (x24 & (x25 | x26)))) | (~x25 & ((~x02 & x23) | (~x22 & ~x24))) | (x23 & (~x24 | (~x02 & ~x22))) | (~x02 & ~x22 & (~x24 | (x25 & x26))))) | (~x22 & ((~x02 & ((x21 & x24 & x25) | (x23 & (x24 | (x25 & x26))))) | (x21 & ((x02 & (~x24 | ~x26)) | (~x23 & ((~x24 & ~x26) | (x02 & x25))))))) | (x21 & ~x23 & ~x24 & ((x22 & ~x25) | (~x02 & ~x26))))) | x04 | (~x11 & x12 & ~x14) | (~x13 & x15) | (x13 & ~x15);
endmodule