module pla__bc0 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10;
  assign z00 = x02 ? (x01 ? (x00 ? ~x03 : (x14 & x15 & (x03 | (~x03 & x04)))) : ((x03 & ((x12 & ((~x00 & x13) | (x00 & x04 & x14 & x15))) | (~x00 & ((x13 & (~x15 | (~x12 & x14 & x15))) | ~x14 | (~x13 & (x15 | (x14 & ~x15))))) | (x00 & (~x04 | (x04 & ~x12 & (~x13 | ~x15 | (x13 & x15))))))) | (x00 & ~x03 & ~x04 & ~x16 & (x13 ? x15 : (~x14 & (x15 | (~x12 & ~x15))))))) : (x03 & ((~x01 & ~x04 & (x00 ? ((~x13 & (x12 | (~x12 & x14 & ~x15))) | (x12 & (x14 | x15)) | (~x12 & ((x15 & ~x16 & (~x05 | ~x06 | ~x07)) | x13 | ~x14))) : ((~x14 ^ x15) & (x12 | x13)))) | (~x00 & x04)));
  assign z01 = (~x01 & ((x03 & (x00 ? (x02 ? (~x04 | (x04 & ~x10 & ((x15 & (x12 ? x14 : x13)) | (~x12 & (~x13 | ~x15))))) : ((~x16 & ((~x05 & ((x04 & x06 & ~x07 & x08 & ~x09 & x10) | (~x04 & ~x12 & x15))) | (~x04 & ~x12 & x15 & (~x06 | ~x07)))) | (~x04 & ((x13 & (~x12 | (x12 & ~x14 & ~x15))) | (~x12 & (~x14 | (~x13 & x14 & ~x15))))))) : (~x10 & (x02 ? ((~x13 & (x15 | (x14 & ~x15))) | ~x14 | (x13 & (x12 | ~x15 | (~x12 & x14 & x15)))) : (~x04 & (~x14 ^ x15) & (x12 | x13)))))) | (x00 & ~x03 & (x02 ? (~x04 & ~x10 & ~x16 & (x13 ? x15 : (~x14 & (x15 | (~x12 & ~x15))))) : ((x11 & (x04 ? (x13 | (x14 & x15)) : (x12 & (x13 | x14)))) | (~x04 & ~x11 & x13 & ~x16 & ((~x12 & x14 & ~x15) | (~x14 & x15)))))))) | (~x00 & ((x01 & (x02 ? (~x10 & x14 & x15 & (x03 | (~x03 & x04))) : (~x03 & ~x04))) | (~x02 & x03 & x04)));
  assign z02 = x02 ? (x00 ? (x01 ? ~x03 : (x03 ? (x04 & ((((x15 & (x12 ? x14 : x13)) | (~x12 & (~x13 | ~x15))) & (x11 | (~x10 & ~x11 & ~x18))) | (x12 & x20 & (~x14 | ~x15)))) : (~x04 & ((~x16 & (x13 ? (x15 ? (x11 | (~x10 & ~x11 & ~x18)) : x20) : ((x15 | (~x12 & ~x15)) & (x14 ? x20 : (x11 | (~x10 & ~x11 & ~x18)))))) | (x16 & (~x12 | x13 | x15)) | (~x15 & x20 & x12 & ~x13))))) : ((x14 & (x03 ? ((x15 & (x01 ? (x11 | (~x10 & ~x11 & ~x19)) : (~x12 & x13 & (x11 | (~x10 & ~x11 & ~x18))))) | (~x01 & ~x13 & ~x15 & (x11 | (~x10 & ~x11 & ~x18)))) : (x04 & x15 & ((x01 & (x11 | (~x10 & ~x11 & ~x19))) | (~x01 & ~x12 & x13 & x20))))) | (x20 & (((~x14 | ~x15) & (x03 ? x01 : x04)) | (~x01 & ~x03 & (~x04 | (x04 & (x12 | ~x13)))))) | (~x01 & x03 & (x11 | (~x10 & ~x11 & ~x18)) & ((x13 & (x12 | ~x15)) | ~x14 | (~x13 & x15))))) : ((~x01 & (x00 ? (x03 ? (x04 ? ((~x16 & ((x20 & ((((x05 & ~x06) | (~x05 & x06 & ~x07 & x08 & x09 & x10)) & (~x11 | ~x12)) | (x11 & x12 & ((~x05 & x06 & ~x07 & x08 & x09 & x10 & (x13 ^ x14)) | (x05 & ~x06 & x13 & x14 & x15))) | (x05 & ~x06 & (~x13 | ~x14)))) | (x05 & ((x06 & ~x07) | (~x06 & x11 & x12 & x13 & x14 & ~x15))) | (~x05 & (x06 ? (~x07 & (~x08 | (x08 & (~x10 | (x10 & (~x09 | (x09 & x11 & x12 & (x13 ^ ~x14)))))))) : x07)))) | (x06 & (x07 | (~x07 & x16))) | (~x06 & ((x16 & (x05 | x07)) | (~x05 & ~x07 & x20)))) : (x12 ? (~x13 | x14 | x15) : ((x15 & ((~x16 & (~x05 | ~x06 | ~x07)) | (~x13 & x14 & (x16 | (x05 & x06 & x07 & ~x16))))) | x13 | ~x14 | (~x13 & x14 & ~x15)))) : (x04 ? (~x11 & x20 & (x12 | (~x12 & (~x14 | x15 | (x14 & ~x15))))) : (x11 ? ((~x14 & ~x15 & x12 & ~x13) | (~x12 & x20)) : ((x20 & ((x12 & ((x13 & ~x15) | (x14 & x15 & ~x16))) | (~x12 & x14 & (~x13 | (x13 & x15 & ~x16))) | (~x14 & (~x13 | ~x15)))) | (x16 & ((x13 & (x15 | (~x12 & x14))) | (x12 & ~x13 & x14))))))) : (x03 & ~x04 & ((x20 & ((x12 & (~x14 ^ ~x15)) | (x13 & x14 & ~x15) | (~x12 & (~x13 | (x13 & ~x14 & x15))))) | ((~x14 ^ x15) & (x12 | x13) & (x11 | (~x10 & ~x11 & ~x18))))))) | (x01 & x20 & (x00 ? (x03 ? x04 : (~x04 | (x04 & (~x13 | (x13 & x14 & ~x15))))) : (x03 ^ x04))) | (~x00 & x03 & x04));
  assign z03 = (~x01 & (x00 ? (x02 ? (x03 ? ((x04 & (((x10 | (~x10 & x11)) & (x12 ? (x14 & x15) : (~x15 | (x13 & x15)))) | (x12 & x20 & (~x14 | ~x15)) | (x10 & ~x12 & ~x13))) | (~x10 & (x12 ? ~x04 : ((~x04 & (x13 | (~x11 & ~x13))) | (x11 & ~x13)))) | (~x04 & x10)) : (x04 ? (~x05 | ~x06 | ~x07 | (x05 & x06 & x07)) : ((x16 & (~x12 | x13 | x15)) | (~x15 & x20 & x12 & ~x13) | (~x16 & ((((x13 & x15) | (~x14 & ~x15 & ~x12 & ~x13)) & (x10 | (~x10 & x11))) | (~x13 & ((x14 & x20 & (x15 | (~x12 & ~x15))) | (x11 & ~x14 & x15))) | (x13 & ~x15 & x20)))))) : (x03 ? (x04 ? ((~x16 & ((x20 & ((((x05 & ~x06) | (~x05 & x06 & ~x07 & x08 & x09 & x10)) & (~x11 | ~x12)) | (x11 & x12 & ((~x05 & x06 & ~x07 & x08 & x09 & x10 & (x13 ^ x14)) | (x05 & ~x06 & x13 & x14 & x15))) | (x05 & ~x06 & (~x13 | ~x14)))) | (~x05 & (x06 ? (~x07 & x08 & (~x10 | (~x09 & x10))) : x07)) | (x05 & ~x06 & x11 & x14 & ~x15 & x12 & x13))) | (x05 & (x06 ? x07 : x16)) | (~x06 & ((~x05 & ~x07 & x20) | (x07 & x16))) | (x06 & ~x07 & x16)) : ((x13 & (x12 ? (~x14 & ~x15) : x11)) | (x12 & (~x13 | x14 | x15)) | (~x12 & ((x15 & ((~x13 & x14 & (x16 | (x05 & x06 & x07 & ~x16))) | (x11 & ~x16 & (~x05 | ~x06 | ~x07)))) | (x11 & (~x14 | (~x13 & x14 & ~x15))))))) : (x04 ? (x11 ? (x13 | (x14 & x15) | (~x13 & (~x14 ^ ~x15))) : (x20 & (x12 | (~x12 & (~x14 | x15 | (x14 & ~x15)))))) : (x11 ? (x12 ? (x13 | x14 | (~x13 & ~x14 & x15)) : x20) : ((x14 & (x12 ? ((~x13 & x16) | (x15 & ~x16 & x20)) : (x13 ? (x16 | (~x16 & (~x15 | (x15 & x20)))) : x20))) | (x13 & ((x15 & (x16 | (~x14 & ~x16))) | (x12 & ~x15 & x20))) | (~x14 & x20 & (~x13 | ~x15))))))) : (x02 ? (x03 ? (((~x13 & (x15 | (x14 & ~x15))) | ~x14 | (x13 & (x12 | ~x15 | (~x12 & x14 & x15)))) & (x11 | (x10 & ~x11))) : (x20 & (~x04 | (x04 & (x12 | ~x13 | (x14 & x15 & ~x12 & x13)))))) : (~x03 | (x03 & ~x04 & ((x20 & ((x12 & (~x14 ^ ~x15)) | (x13 & x14 & ~x15) | (~x12 & (~x13 | (x13 & ~x14 & x15))))) | ((~x14 ^ x15) & (x12 | x13) & (x10 | (~x10 & x11))))))))) | (x01 & (x00 ? (x02 | (~x02 & (x03 ? (x04 & x20) : (x04 ? (x13 ? (x14 & (x15 | (~x15 & x20))) : x20) : x20)))) : ((x20 & ((x03 & (x02 ? (~x14 | ~x15) : ~x04)) | (~x02 & ~x03 & x04))) | (x02 & ((~x03 & ~x04) | (x14 & x15 & (x03 ? (x11 | (x10 & ~x11)) : (x04 & (x10 | (~x10 & x11)))))))))) | (~x00 & x04 & (x02 ? (~x03 & x20 & (~x14 | ~x15)) : (x03 & x10)));
  assign z04 = (~x04 & ((~x03 & (x00 ? (~x01 & ~x02 & (x11 ? (x12 & (x13 | x14 | (~x13 & ~x14 & ~x15))) : (~x16 & ((x13 & ~x14 & x15) | (x14 & ~x15 & x12 & ~x13))))) : (x01 | (~x01 & ~x02)))) | (x00 & ~x01 & x03 & (x02 | (~x02 & x12 & (~x13 | x14 | x15 | (x13 & ~x14 & ~x15))))))) | (x00 & ((~x03 & ((x02 & (x01 | (x05 & x06 & x07 & ~x01 & x04))) | (~x01 & ~x02 & x04 & x11 & (x13 | (x14 & x15))))) | (~x01 & ~x02 & x03 & x04 & ((~x16 & (x05 ? ((x06 & ~x07) | (~x06 & x11 & x12 & x13 & x14 & ~x15)) : (x06 ? (~x07 & x08 & (x09 ? (~x10 | (x10 & x11 & x12 & x13 & x14)) : x10)) : x07))) | (~x05 & x06 & x07)))));
  assign z05 = (~x02 & ((~x03 & (x00 ? ((~x01 & (x04 ? (x11 & (x13 | (x14 & x15) | (~x13 & ((~x14 & x15) | (x12 & x14 & ~x15))))) : (x11 ? (x12 & (x13 | x14 | (~x13 & ~x14 & x15))) : (~x16 & ((x13 & ~x14 & x15) | (x14 & ~x15 & x12 & ~x13)))))) | (x13 & x15 & x01 & x04)) : (x01 ^ x04))) | (x00 & x03 & ((~x09 & ((x01 & ~x04 & ~x08 & ~x10) | (~x01 & x04 & ~x05 & x06 & ~x07 & x08 & x10 & ~x15 & ~x16))) | (~x01 & x04 & ((~x05 & x06 & x07) | (~x16 & ((x05 & ~x06 & x11 & x14 & ~x15 & x12 & x13) | (~x05 & (x06 ? (~x07 & x08 & (~x10 | (x12 & x13 & x14 & x09 & x10 & x11))) : x07)))))) | (x01 & ~x04 & (((~x14 | x15) & (x08 | x09 | x10) & (x05 | x06 | x07)) | (x14 & ~x15) | (~x05 & ~x06 & ~x07))))))) | (x01 & x02 & (x00 ? x03 : (~x10 & ~x11 & x14 & x15 & ~x19 & (x03 | (~x03 & x04)))));
  assign z06 = (~x01 & (x00 ? (x03 ? (x02 ? (~x04 | (x04 & ((x15 & (x12 ? x14 : x13)) | (~x12 & (~x13 | ~x15))))) : ((~x16 & ((~x06 & (x04 ? (~x05 & x07) : (~x12 & x15))) | (x15 & ((~x04 & ~x12 & (~x05 | ~x07)) | (x06 & ~x07 & x04 & ~x05 & x08 & ~x09 & x10 & x11 & ~x13))) | (x04 & ~x05 & x06 & ~x07 & x08 & (~x10 | (x10 & x11 & ~x14 & (x09 ? (x12 & ~x13) : ~x15)))))) | (~x04 & ((x13 & (~x12 | (x12 & ~x14 & ~x15))) | (~x12 & (~x14 | (~x13 & x14 & ~x15))) | (x12 & (~x13 | x14 | x15)))) | (x06 & x07 & x04 & ~x05))) : (x04 ? ((x02 & (~x05 | ~x06 | ~x07 | (x05 & x06 & x07))) | (~x13 & ~x14 & ~x15 & ~x02 & x11)) : (~x16 & ((x13 & (x02 ? x15 : (~x11 & ((~x12 & x14 & ~x15) | (~x14 & x15))))) | (x02 & ~x13 & ~x14 & (x15 | (~x12 & ~x15))))))) : (x03 & (x02 ? ((~x13 & (x15 | (x14 & ~x15))) | ~x14 | (x13 & (x12 | ~x15 | (~x12 & x14 & x15)))) : (~x04 & (~x14 ^ x15) & (x12 | x13)))))) | (~x00 & ((x01 & x02 & x14 & x15 & (x03 | (~x03 & x04))) | (~x02 & (x03 ^ ~x04)))) | (x00 & x01 & ~x03 & (x02 | (~x02 & x04 & x13 & (x15 | (~x14 & ~x15)))));
  assign z07 = x00 ? (x02 ? (x01 | (~x01 & (x03 ? (~x04 | (x04 & x12 & ((x14 & x15) | (x20 & (~x14 | ~x15))))) : (x04 ? (~x05 | ~x06 | ~x07) : ((x16 & (~x12 | x13 | x15)) | (~x15 & x20 & x12 & ~x13) | (~x16 & (x13 ? (x15 ? ~x12 : x20) : ((x15 | (~x12 & ~x15)) & (~x14 | (x14 & x20)))))))))) : (x03 ? ((~x08 & ((x01 & ~x04 & ~x09 & ~x10) | (~x01 & x04 & ~x05 & x06 & ~x07 & ~x16))) | (~x01 & (x04 ? ((x07 & (x06 ? x05 : x16)) | (~x16 & (x05 ? (~x06 & x20 & (~x11 | ~x12 | ~x13 | ~x14 | (x11 & x12 & x13 & x14 & x15))) : (x06 & ~x07 & x08 & (~x10 | (x10 & (((x13 ^ x14) & ((~x09 & x15) | (x09 & x11 & x12 & x20))) | (x09 & ((x11 & x12) ? (x13 & x14 & x15) : x20)))))))) | (x06 & ~x07 & x16) | (~x06 & (x05 ? x16 : (~x07 & x20)))) : ((~x15 & (x12 ? (x13 & ~x14) : (~x13 & x14))) | (x12 & (x14 | x15)) | (~x13 & (x12 | (~x12 & x14 & x15 & (x16 | (x05 & x06 & x07 & ~x16)))))))) | (x01 & (x04 ? x20 : (((~x14 | x15) & (x08 | x09 | x10) & (x05 | x06 | x07)) | (x14 & ~x15) | (~x05 & ~x06 & ~x07))))) : ((x20 & (x01 ? (~x04 | (x04 & (~x13 | (x13 & x14 & ~x15)))) : ((~x11 & (x04 ? (x12 | (~x12 & (~x14 | x15 | (x14 & ~x15)))) : ((x12 & ((x13 & ~x15) | (x14 & x15 & ~x16))) | (~x12 & x14 & (~x13 | (x13 & x15 & ~x16))) | (~x14 & (~x13 | ~x15))))) | (~x04 & x11 & ~x12)))) | (~x01 & ((~x13 & ((x14 & ((~x04 & ~x11 & x12 & (x16 | (~x15 & ~x16))) | (~x12 & ~x15 & x04 & x11))) | (x04 & x11 & ~x14 & (~x15 | (~x12 & x15))))) | (~x04 & ~x11 & x13 & x16 & (x15 | (~x12 & x14)))))))) : ((x20 & ((~x01 & ((~x13 & ((x02 & ~x03 & x04) | (~x02 & x03 & ~x04 & ~x12))) | (x02 & ~x03 & (~x04 | (x04 & (x12 | (x14 & x15 & ~x12 & x13))))) | (~x02 & x03 & ~x04 & ((x12 & (~x14 ^ ~x15)) | (x13 & ((x14 & ~x15) | (~x12 & ~x14 & x15))))))) | (x01 & ((x03 & (x02 ? (~x14 | ~x15) : ~x04)) | (~x02 & ~x03 & x04))) | (x02 & ~x03 & x04 & (~x14 | ~x15)))) | (~x01 & ((~x02 & ~x03 & ~x04) | (x13 & x14 & x15 & x02 & x03 & ~x12))) | (x01 & ((x03 & (x02 ? (x14 & x15) : x04)) | (x02 & ~x03 & (~x04 | (x04 & x14 & x15))))));
  assign z08 = x00 ? ((~x02 & (x03 ? ((~x10 & ((x01 & ~x04 & ~x08 & ~x09) | (~x01 & x04 & ~x05 & x06 & ~x07 & x08 & x09 & ~x16))) | (x01 & (x04 ? x20 : (((~x14 | x15) & (x08 | x09 | x10) & (x05 | x06 | x07)) | (x14 & ~x15) | (~x05 & ~x06 & ~x07)))) | (~x01 & (x04 ? (x06 ? (~x07 & (x16 | (~x16 & (x05 | (~x05 & x08 & x09 & x10 & x20 & (~x11 | ~x12 | (x11 & x12 & (x13 ^ x14)))))))) : ((x07 & (x16 | (x05 & x11 & x12 & x13 & x14 & ~x15 & ~x16))) | (~x05 & ~x07 & x20) | (x05 & (x16 | (~x16 & x20 & (~x11 | ~x12 | ~x13 | ~x14 | (x11 & x12 & x13 & x14 & x15))))))) : ((x13 & (~x12 | (~x14 & ~x15 & x11 & x12))) | (x12 & ~x17 & (~x13 | x14 | x15)) | (~x12 & ((~x13 & x14 & (~x15 | (x15 & x16))) | ~x14 | (x15 & ~x16 & (~x05 | ~x06 | ~x07)))))))) : (x01 ? (x04 ? (x13 ? (x15 | (~x15 & (~x14 | (x14 & x20)))) : x20) : x20) : (x11 ? ((~x13 & (x04 ? (x12 ? (x14 & ~x15) : ~x14) : (x12 & ~x14))) | (~x04 & ~x12 & x20)) : ((x20 & (x04 ? (x12 | (~x12 & (~x14 | x15 | (x14 & ~x15)))) : ((x12 & ((x13 & ~x15) | (x14 & x15 & ~x16))) | (~x12 & x14 & (~x13 | (x13 & x15 & ~x16))) | (~x14 & (~x13 | ~x15))))) | (~x04 & x16 & ((x13 & (x15 | (~x12 & x14))) | (x12 & ~x13 & x14)))))))) | (~x01 & x02 & ((~x14 & ((~x03 & ~x04 & ~x12 & ~x13 & ~x15 & ~x16) | (x03 & x04 & x12 & x20))) | (x04 & (x03 ? (x12 ? (x15 ? x14 : x20) : (~x13 | ~x15 | (x13 & x15))) : (~x05 | ~x06 | ~x07 | (x05 & x06 & x07)))) | (~x04 & (x03 ? x13 : ((~x12 & (x16 | (~x13 & x14 & ~x15 & ~x16 & x20))) | (x20 & (x13 ? (~x15 & ~x16) : ((x14 & x15 & ~x16) | (x12 & ~x15)))) | (x15 & x16) | (x13 & (x16 | (x15 & ~x16))))))))) : ((~x01 & (x02 ? ((x12 & (x03 ? x13 : (x04 & x20))) | (~x03 & x20 & (~x04 | (x04 & (~x13 | (x14 & x15 & ~x12 & x13))))) | (x03 & ((x13 & (~x15 | (~x12 & x14 & x15))) | ~x14 | (~x13 & (x15 | (x14 & ~x15)))))) : (x03 ? (~x04 & (((~x14 ^ x15) & (x12 | x13)) | (x20 & ((x12 & (~x14 ^ ~x15)) | (x13 & x14 & ~x15) | (~x12 & (~x13 | (x13 & ~x14 & x15))))))) : x04))) | (x01 & ((x20 & ((x03 & (x02 ? (~x14 | ~x15) : ~x04)) | (~x02 & ~x03 & x04))) | (x02 & x14 & x15 & (x03 | (~x03 & x04))))) | (x04 & (x02 ? (~x03 & x20 & (~x14 | ~x15)) : x03)));
  assign z09 = x03 ? (x02 ? (x00 ? (~x01 & (x04 ? (~x12 & (~x13 | ~x15 | (x13 & x15))) : ~x14)) : ((~x01 & (~x14 | (~x13 & (x15 | (x14 & ~x15))) | (x13 & (x12 | ~x15)))) | (x01 & ~x10 & ~x11 & x14 & x15))) : (x00 ? ((~x08 & ((~x01 & x04 & ~x05 & x06 & ~x07 & ~x16) | (x01 & ~x04 & ~x09 & ~x10 & ~x12))) | (~x01 & ((~x16 & ((x06 & ((x05 & ((x04 & ~x07) | (~x04 & x07 & ~x12 & ~x13 & x14 & x15))) | (x04 & ~x05 & ~x07 & x08 & x10 & (~x09 | (x09 & x11 & x12 & (x13 ? x14 : (~x14 & ~x15))))))) | (~x04 & ~x12 & x15 & (~x06 | ~x07)) | (~x05 & (x04 ? (~x06 & x07) : (~x12 & x15))))) | (~x04 & (x12 ? ((~x17 & (~x13 | x14 | x15)) | (~x14 & ~x15 & ~x11 & x13)) : (x13 | ~x14))))) | (x01 & ~x04 & ~x12 & (((~x14 | x15) & (x08 | x09 | x10) & (x05 | x06 | x07)) | (x14 & ~x15) | (~x05 & ~x06 & ~x07)))) : (~x01 & (x04 | (~x04 & (~x14 ^ x15) & (x12 | x13)))))) : ((x01 & (x00 ? (x02 | (~x02 & x04 & x13 & (x15 | (~x14 & ~x15)))) : ((~x02 & ~x04) | (~x11 & x14 & x15 & x02 & x04 & ~x10)))) | (x00 & ~x01 & ((~x02 & ((x11 & ~x13 & ((x04 & (x15 ? ~x14 : ~x12)) | (~x14 & ~x15 & ~x04 & x12))) | (x13 & x14 & ~x15 & ~x16 & ~x04 & ~x11 & ~x12))) | (x13 & x15 & ~x16 & x02 & ~x04 & x12))));
  assign z10 = (~x01 & (x00 ? (x02 ? ((x20 & ((x12 & ((x03 & x04 & (~x14 | ~x15)) | (~x03 & ~x04 & ~x13 & ~x15))) | (~x03 & ~x04 & ~x16 & (x13 ? ~x15 : (x14 & (x15 | (~x12 & ~x15))))))) | (x03 & ~x04 & x15)) : (x03 ? (x04 ? ((x07 & (x05 ? x06 : (~x06 & ~x16))) | (~x16 & ((x06 & ~x07 & (x05 | (~x05 & (~x08 | (x08 & (x09 ? (~x10 | (x10 & ((x20 & (~x11 | ~x12)) | (x11 & x12 & (x13 ? (x14 | (~x14 & x20)) : (x14 & x20)))))) : (x10 ? x14 : x15))))))) | (x05 & ~x06 & ((x11 & x12 & x13 & x14 & (~x15 | (x15 & x20))) | (x20 & (~x11 | ~x12 | ~x13 | ~x14)))))) | (~x07 & x20 & ~x05 & ~x06)) : ((~x13 & ((x11 & x12) | (x05 & x06 & x07 & x15 & ~x16 & ~x12 & x14))) | (x11 & x12 & (x14 | x15 | (x13 & ~x14 & ~x15))))) : ((~x12 & (x11 ? ((~x04 & x20) | (~x14 & x15 & x04 & ~x13)) : (x20 & ((x14 & (x04 ? ~x15 : (~x13 | (x13 & x15 & ~x16)))) | (x04 & (~x14 | x15)))))) | (~x11 & (x04 ? (x12 & x20) : ((x13 & ((x12 & ~x15 & x20) | (~x14 & x15 & ~x16))) | (~x14 & x20 & (~x13 | ~x15)) | (x12 & x14 & ~x16 & (x15 ? x20 : ~x13))))) | (x11 & x12 & ~x13 & ~x14 & ~x15)))) : ((~x02 & ~x03 & ~x04) | (x20 & ((~x13 & ((x02 & ~x03 & x04) | (~x02 & x03 & ~x04 & ~x12))) | (x02 & ~x03 & (~x04 | (x04 & (x12 | (x14 & x15 & ~x12 & x13))))) | (~x02 & x03 & ~x04 & ((x12 & (~x14 ^ ~x15)) | (x13 & ((x14 & ~x15) | (~x12 & ~x14 & x15)))))))))) | (x01 & (x02 ? (x00 ? ~x03 : (x03 & x20 & (~x14 | ~x15))) : ((x20 & (x00 ? (x03 ? x04 : (~x04 | (x04 & (~x13 | (x13 & x14 & ~x15))))) : (x03 ^ x04))) | (x00 & ~x03 & x04 & x13 & (x15 | (~x14 & ~x15)))))) | (~x00 & x02 & ~x03 & x04 & x20 & (~x14 | ~x15));
endmodule