module pla__mp2d ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13;
  assign z00 = ~x00 | (x00 & (x01 | (~x01 & (~x02 | (x02 & (x03 | (~x03 & (~x04 | (x04 & (~x05 | (x05 & (x06 | (~x06 & (~x07 | (x07 & (x08 | (~x08 & (x09 | (~x09 & x10)))))))))))))))))));
  assign z01 = ((x06 | (~x06 & (~x07 | (x07 & (x08 | (~x08 & (x09 | (~x09 & ~x10)))))))) & (~x00 | (x00 & ((x01 & (x02 | (~x02 & ~x03 & ~x04))) | (~x01 & ~x03 & (x02 | (~x02 & x04))) | (~x02 & x03))))) | (x00 & ((~x01 & (x02 ? x03 : (~x03 & ~x04))) | (x01 & ~x02 & ~x03 & x04)));
  assign z02 = (x00 & ((~x03 & (x01 ? (~x05 | (~x02 & (x04 | (~x04 & (x06 | (~x06 & (~x07 | (x07 & (x08 | (~x08 & (~x09 | (x09 & x10)))))))))))) : ((~x04 & (~x02 | (x02 & ~x05))) | ((x02 | (~x02 & x04)) & (x06 | (~x06 & (~x07 | (x07 & (x08 | (~x08 & (~x09 | (x09 & x10))))))))) | (x02 & x04) | (~x02 & ~x05)))) | (x01 & x02 & (x06 | (~x06 & (~x07 | (x07 & (x08 | (~x08 & (~x09 | (x09 & x10))))))))))) | x03 | (~x00 & ((~x06 & (~x07 | (x07 & (x08 | (~x08 & (~x09 | (x09 & x10))))))) | x06 | (~x03 & ~x05)));
  assign z03 = (x00 & ((~x01 & (x02 ? x03 : (~x03 & ~x04))) | (x01 & ~x02 & ~x03 & x04))) | ((~x00 | (x00 & ((x01 & (x02 | (~x02 & ~x03 & ~x04))) | (~x01 & ~x03 & (x02 | (~x02 & x04))) | (~x02 & x03)))) & (x06 | (~x06 & (~x07 | (x07 & (x08 | (~x08 & (~x09 | (x09 & ~x10)))))))));
  assign z04 = (x00 & ((~x01 & ((x02 & x03) | (~x02 & ~x03 & ~x04 & x08 & ~x09 & ~x10))) | (x01 & ~x02 & ~x03 & ~x09 & ~x10 & x04 & x08))) | (x08 & ~x09 & ~x10 & (x06 | (~x06 & ~x07)));
  assign z05 = (x00 & ((~x01 & (x02 ? x03 : (~x03 & ~x04))) | (x01 & ~x02 & ~x03 & x04))) | ((~x00 | (x00 & ((x01 & (x02 | (~x02 & ~x03 & ~x04))) | (~x01 & ~x03 & (x02 | (~x02 & x04))) | (~x02 & x03)))) & (x06 | (~x06 & (~x07 | (x07 & (~x08 | (x08 & (x09 | (~x09 & ~x10)))))))));
  assign z06 = x00 & x07 & ((~x01 & (x02 ? x03 : (~x03 & ~x04))) | (x01 & ~x02 & ~x03 & x04)) & (~x06 | (x09 & x10 & x06 & x08));
  assign z07 = ~x04 & ~x03 & ~x02 & x00 & ~x01;
  assign z08 = x04 & ~x03 & ~x02 & x00 & x01;
  assign z09 = (x00 & ((~x01 & (x02 ? x03 : (~x03 & ~x04))) | (x01 & ~x02 & ~x03 & x04))) | ~x06 | (x06 & (~x07 | (x07 & (~x08 | (x08 & (~x09 | (x09 & ~x10)))))));
  assign z10 = (~x00 & ~x01 & ((~x03 & x04) | (x02 & x03 & ~x04))) | (x00 & x01 & ~x02 & ~x03 & x04);
  assign z11 = ~x13 & x12 & ~x11 & x10 & x09 & x08 & x06 & x07;
  assign z12 = ~x13 & x12 & ~x11 & x10 & x09 & x08 & x06 & x07;
  assign z13 = x00 | (~x00 & (~x01 | (x01 & (~x02 | (x02 & (~x03 | (x03 & x04)))))));
endmodule