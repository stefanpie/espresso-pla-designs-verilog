module pla__jbp ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56;
  assign z00 = x20 & ~x29 & ~x30 & ~x34 & (x00 | (x08 & (~x01 | x09)));
  assign z01 = (~x00 & x01 & ~x09 & x20 & ~x29 & ~x30 & ~x34 & (x08 | (x03 & x10 & x11 & ~x12 & ~x13))) | (x28 & x29);
  assign z02 = (~x00 & x20 & ~x29 & ~x30 & ~x34 & ((x09 & (x01 | ~x08)) | (x01 & ~x08 & ~x13 & (x10 ? (~x03 | (x11 & ~x12)) : (~x11 & ~x12))))) | (~x28 & x29);
  assign z03 = (~x32 & ((~x26 & ((~x27 & ((~x21 & x28 & (x22 ? (~x29 & ~x33) : (x23 ? (~x29 & x33) : (x29 & (x24 ^ x33))))) | (x21 & ~x28 & x29 & x33))) | (x27 & ~x28 & x29 & ~x33))) | (~x29 & x33 & x26 & ~x28))) | ~x31 | (~x28 & ~x29 & x32 & ~x33);
  assign z04 = x16 & x25;
  assign z05 = ~x34 & ~x30 & ~x29 & x20 & ~x13 & x12 & x10 & ~x09 & ~x08 & ~x03 & ~x00 & x01;
  assign z06 = x00 & ~x29 & ~x30 & ((x09 & ((~x01 & ((x08 & ~x10 & x11 & x12) | (~x11 & x13))) | (x12 & x13))) | (x10 & x13));
  assign z07 = ~x29 & ~x30 & ((x00 & x01 & ~x13 & (x10 | (x09 & (~x11 | x12)))) | (~x09 & ~x10 & x12 & (x08 | ~x11)));
  assign z08 = x29 | (~x30 & ((x09 & (x01 ? (~x10 & ~x11 & x13 & (x00 | ~x12)) : (~x13 & ((x08 & ~x10 & x11 & x12) | (~x00 & (~x11 | x12)))))) | (~x08 & ~x09 & ~x10 & x11 & x12) | (~x00 & ~x01 & x10 & ~x13)));
  assign z09 = ~x29 & ((~x00 & (~x01 | (x12 & x13))) | (~x10 & (~x09 | (x11 & ~x12))) | x30 | (x13 & (~x01 | x10 | x11)));
  assign z10 = x29 | (~x30 & ((x12 & ((x09 & (x00 ? ((~x08 & x11) | (x01 & ~x13)) : (~x01 & x13))) | (~x10 & ((x08 & (~x09 | (~x00 & ~x01 & x11))) | (~x09 & ~x11))))) | (~x01 & ((x10 & x13) | (x00 & x09 & ~x11))) | (x00 & (x10 | (x09 & ~x11 & ~x12))) | (x09 & ~x10 & ~x11 & ~x12 & x13)));
  assign z11 = ~x29 & ~x30 & (x10 | (x09 & (~x11 | x12)));
  assign z12 = (x07 & ~x11 & x30) | (~x00 & x01 & x03 & ~x08 & ~x09 & ~x10 & x11 & x12 & ~x13 & x20 & ~x29 & ~x30 & ~x34);
  assign z13 = ~x34 & ~x30 & ~x29 & x20 & x09 & ~x08 & ~x00 & x01;
  assign z14 = ~x00 & x01 & ~x08 & ~x09 & ~x13 & x20 & ~x29 & ~x30 & ~x34 & (x10 ? (x03 ? x11 : x12) : (~x11 & x12));
  assign z15 = x29 & x19 & x28;
  assign z16 = x34 & ~x30 & ~x28 & ~x29;
  assign z17 = ~x34 & ~x30 & ~x29 & x20 & ~x09 & x08 & ~x00 & x01;
  assign z18 = (x07 & ~x11 & x30) | (x11 & ((~x07 & x30) | (~x00 & x01 & x03 & ~x08 & ~x09 & ~x10 & ~x13 & x20 & ~x29 & ~x30 & ~x34)));
  assign z19 = (~x28 & x29) | (~x00 & ~x01 & x08 & x13 & x14 & x15 & (x29 | (x20 & ~x30 & ~x34)) & (x02 ^ x03));
  assign z20 = x31;
  assign z21 = ~x16 & x25;
  assign z22 = x01 ? x08 : ((~x08 & ((x03 & x07 & ~x09) | (~x11 & ~x12 & x09 & ~x10))) | (~x10 & ~x11 & ~x12 & ~x07 & x09));
  assign z23 = (x07 & (x01 | (~x08 & ((~x11 & ~x12 & x09 & ~x10) | (x04 & ~x09))))) | (~x10 & ~x11 & x12 & ~x01 & ~x07 & x09);
  assign z24 = (x07 & ~x08 & ((~x11 & ~x12 & x09 & ~x10) | (~x01 & x05 & ~x09))) | (x09 & (x01 | (x11 & ~x12 & ~x07 & ~x10)));
  assign z25 = x01 ? x13 : ((x07 & ~x08 & ((~x11 & ~x12 & x09 & ~x10) | (x06 & ~x09))) | (~x10 & x11 & x12 & ~x07 & x09));
  assign z26 = x01 ? x14 : ((x07 & ~x08 & ((x03 & x09) | (~x11 & ~x12 & ~x09 & ~x10))) | (~x07 & x09 & x10 & ~x11 & ~x12));
  assign z27 = x01 ? x15 : ((x07 & ~x08 & ((~x11 & ~x12 & ~x09 & ~x10) | (x04 & x09))) | (~x07 & x09 & x10 & ~x11 & x12));
  assign z28 = x01 ? x00 : ((x07 & ~x08 & ((~x11 & ~x12 & ~x09 & ~x10) | (x05 & x09))) | (~x07 & x09 & x10 & x11 & ~x12));
  assign z29 = x01 ? x02 : ((x07 & ~x08 & ((~x11 & ~x12 & ~x09 & ~x10) | (x06 & x09))) | (~x07 & x09 & x10 & x11 & x12));
  assign z30 = x30 | (~x00 & x01 & x03 & ~x08 & ~x09 & x11 & ~x13 & x20 & ~x29 & ~x34 & (~x10 | x12));
  assign z31 = (~x28 & x29) | (~x00 & x01 & ~x08 & ~x09 & x10 & ~x13 & x20 & ~x29 & ~x30 & ~x34 & (~x03 | (x11 & ~x12)));
  assign z32 = ~x31 | (~x21 & ~x26 & ~x27 & ~x32);
  assign z33 = ~x32 & x31 & ~x27 & ~x21 & ~x26;
  assign z34 = ~x31 | (~x26 & ~x32 & (x21 | x27 | (~x22 & ~x23)));
  assign z35 = ~x26 & x31 & ~x32 & (x21 | x27 | (~x22 & ~x23));
  assign z36 = x31 & (x32 | (~x26 & (x27 | (~x21 & (x22 | (~x23 & x24))))));
  assign z37 = x31 & ~x32 & (x26 | (~x27 & (x21 | (~x22 & (x23 | ~x24)))));
  assign z38 = ~x34 & ~x30 & ~x29 & x20 & x09 & ~x00 & ~x08;
  assign z39 = ~x34 & ~x30 & ~x29 & x20 & ~x13 & x10 & ~x09 & ~x08 & ~x03 & ~x00 & x01;
  assign z40 = ~x34 & ~x30 & ~x29 & x20 & ~x13 & ~x11 & ~x10 & ~x09 & ~x08 & x03 & ~x00 & x01;
  assign z41 = x00 & ~x29 & ~x30 & ((x13 & ((x01 & x17 & (x10 | (x09 & x12))) | (~x10 & x11 & x12 & ~x01 & x08 & x09))) | (~x01 & x08 & x09 & ~x10 & x11 & x12 & x17));
  assign z42 = ~x34 & ~x30 & ~x29 & x20 & ~x13 & x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x00 & x01;
  assign z43 = ~x34 & ~x30 & ~x29 & x20 & ~x13 & ~x11 & ~x10 & ~x09 & ~x08 & ~x00 & x01;
  assign z44 = ~x00 & x08 & x09 & x20 & ~x29 & ~x30 & ~x34 & (x01 | (x10 & x11 & ~x12));
  assign z45 = x20 & ~x29 & ~x30 & ~x34 & (x00 | (x01 & x09) | (~x01 & x08 & x10 & x11 & x12));
  assign z46 = ~x00 & x01 & ~x08 & ~x09 & x13 & x20 & ~x29 & ~x30 & ~x34 & ((~x11 & (x10 ? (x12 ^ x18) : (x12 ^ x35))) | (~x10 & x11 & (x12 ^ x17)));
  assign z47 = x20 & ~x29 & ~x30 & ~x34 & (((~x10 | x12) & (x00 | (x01 & x08 & x09))) | (x08 & x10 & x11 & ((x09 & x12) | (~x00 & ~x01 & ~x09 & ~x12))) | (x01 & ~x08 & ~x09 & ~x10 & ~x11 & x12 & ~x13));
  assign z48 = x28 & x29;
  assign z49 = ~x34 & ~x30 & ~x29 & x20 & ~x13 & ~x12 & x10 & ~x09 & ~x08 & ~x03 & ~x00 & x01;
  assign z50 = ~x34 & ~x30 & ~x29 & x20 & ~x13 & ~x12 & ~x11 & ~x10 & ~x09 & ~x08 & ~x00 & x01;
  assign z51 = (x20 & ~x34 & (((~x10 | x12) & (x00 | (x01 & x08))) | (~x09 & ((~x00 & ((x01 & (x08 | (x03 & x11 & ~x13))) | (x11 & ~x12 & x08 & x10))) | (x01 & x12 & ~x13 & (x10 ? ~x03 : ~x11)))) | (x10 & x11 & x12 & x08 & x09))) | x29 | x30;
  assign z52 = ~x00 & ~x01 & x20 & ~x29 & ~x30 & ~x34 & (x08 | x09);
  assign z53 = ~x28 & x29;
  assign z54 = ~x00 & ~x09 & x20 & ~x29 & ~x30 & ~x34 & (~x01 ^ x08);
  assign z55 = ~x00 & ~x01 & x08 & x20 & ~x29 & ~x30 & ~x34 & (~x10 | x12);
  assign z56 = x30 | (~x00 & x01 & x03 & ~x08 & ~x09 & ~x10 & x11 & ~x13 & x20 & ~x29 & ~x34);
endmodule