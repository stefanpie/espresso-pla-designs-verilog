module pla__in6 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22;
  assign z00 = ~x00 & ((~x15 & ~x16 & x31) | (x01 & x22 & x28 & x30 & ~x31));
  assign z01 = ~x00 & ((~x04 & x32) | (x01 & x24 & x28 & x29 & ~x32));
  assign z02 = ~x30 & ~x28 & ~x00 & x03;
  assign z03 = x00 | (~x00 & x03 & ~x28 & x29 & ~x30);
  assign z04 = ~x00 & ~x28 & x30 & ((~x10 & ((~x09 & x11 & ~x12) | (x09 & x19 & x20 & x21 & x29))) | (x10 & (x09 ? (x11 ? (x19 & x29 & (x12 ? x20 : x21)) : x12) : ((~x11 & ~x12) | (x21 & x29 & x11 & x12)))) | (x09 & ~x11 & ~x12 & x21 & x29 & x19 & x20));
  assign z05 = ~x00 & ~x16 & ~x18 & x30 & ((x01 & x23 & x28 & ((~x06 & ((~x15 & x17) | (x07 & x15 & ~x17))) | (~x14 & x15 & x17))) | (~x11 & ~x12 & ~x09 & x10 & ~x14 & x15 & x17 & ~x28));
  assign z06 = ~x00 & ~x15 & x30 & ((((x16 & ~x17 & x18) | (~x06 & ~x16 & x17 & ~x18)) & ((x01 & x23 & x28) | (~x09 & x10 & ~x11 & ~x12 & ~x28))) | (x01 & ~x09 & ~x10 & x11 & x12 & ~x16 & x23 & ~x28 & (x17 ? (x06 | (~x06 & ~x08 & x18)) : ~x18)));
  assign z07 = x00 | (x16 & ~x17 & x30 & ((~x00 & ~x15 & x18 & ((~x09 & x10 & ~x11 & ~x12 & ~x28) | (x01 & x22 & x28))) | (x01 & x15 & ~x18 & x22 & (x28 | (x11 & x12 & ~x09 & ~x10)))));
  assign z08 = x00 | (x15 & ~x18 & x30 & ((~x09 & ~x28 & ((~x00 & ((x10 & ~x11 & ~x12 & ~x14 & ~x16 & x17) | (x01 & ~x06 & x08 & ~x10 & x11 & x12 & x16 & ~x17 & x22))) | (~x06 & x07 & x10 & ~x11 & ~x12 & ~x16 & ~x17))) | (x01 & x22 & x28 & (~x16 | (x16 & ~x17)))));
  assign z09 = (~x16 & ~x18 & x30 & ((x01 & x22 & x28 & ((~x00 & x17 & (x15 ? ~x14 : ~x06)) | (x15 & ~x17 & ~x06 & x07))) | (~x00 & ~x09 & x10 & ~x11 & ~x12 & ~x14 & x15 & x17 & ~x28))) | (x00 & x07);
  assign z10 = (x00 & x07) | (~x17 & x30 & ((x01 & x22 & ((~x18 & ((~x09 & ~x10 & x11 & x12 & ~x28 & ((~x00 & ((x06 & (x15 | ~x16)) | (~x06 & x08 & x15 & x16))) | (x07 & ~x15 & ~x16))) | (~x06 & x07 & x15 & ~x16 & x28))) | (~x00 & ~x15 & x16 & x18 & x28))) | (~x09 & x10 & ~x11 & ~x12 & ~x28 & ((~x00 & ~x15 & x16 & x18) | (~x06 & x07 & x15 & ~x16 & ~x18)))));
  assign z11 = x00 ? ~x07 : (~x15 & x18 & x30 & ((~x09 & ((x01 & ~x10 & x11 & x12 & ~x16 & x17 & x23) | (x10 & ~x11 & ~x12 & x16 & ~x17 & ~x28))) | (x01 & x23 & x28 & (x16 ^ x17))));
  assign z12 = x00 ? ~x07 : (~x16 & x17 & x30 & ((~x09 & ~x28 & ((~x06 & ~x15 & ((x10 & ~x11 & ~x12 & ~x18) | (x01 & ~x08 & ~x10 & x11 & x12 & x18 & x23))) | (x10 & ~x11 & ~x12 & ~x14 & x15 & ~x18))) | (x01 & x23 & x28 & (~x18 | (~x15 & x18)))));
  assign z13 = x00 | (x01 & x28 & x29 & (x25 | (~x00 & x24)));
  assign z14 = x29 & x28 & x24 & ~x22 & x13 & ~x00 & x01;
  assign z15 = x29 & x28 & x24 & ~x00 & x01;
  assign z16 = ~x00 & (x05 | (x22 & x28 & x30));
  assign z17 = (x26 & (~x03 | x27)) | x00 | (~x00 & ~x09 & x10 & ~x11 & ~x12 & ~x28 & x30);
  assign z18 = x00 | (~x03 & x27) | (~x00 & ~x09 & x10 & ~x11 & ~x12 & ~x28 & x30) | (x03 & x26 & ~x27);
  assign z19 = ~x00 & ~x28 & x30 & ((x11 & ((x10 & x29 & (x09 ? (x19 & (x12 ? x20 : x21)) : (x12 & x21))) | (~x09 & ~x10 & ~x12))) | (x09 & ((~x11 & ((x10 & x12) | (x20 & x21 & x29 & ~x12 & x19))) | (x20 & x21 & x29 & ~x10 & x19))));
  assign z20 = x00 | (~x28 & ((~x00 & ((x30 & ((x09 & (x10 ? ((~x11 & x12) | (x11 & ~x12 & x19 & x21 & x29)) : (x19 & x20 & x21 & x29 & (~x12 | (x11 & x12))))) | (~x09 & x10 & x11 & x12 & x21 & x29))) | (x03 & ~x29 & ~x30))) | (~x30 & (x29 ? ~x03 : x02))));
  assign z21 = ~x00 & ~x28 & (x30 ? ((~x10 & ((~x09 & x11 & ~x12) | (x20 & x21 & x29 & x09 & x12 & x19))) | (x09 & x19 & x20 & x29 & ((x10 & x11 & x12) | (~x11 & ~x12 & x21)))) : x03);
  assign z22 = x30 & x29 & ~x28 & x20 & x19 & x12 & x11 & x10 & ~x00 & x09;
endmodule