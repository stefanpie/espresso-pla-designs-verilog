module pla__t3 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11,
    z0, z1, z2, z3, z4, z5, z6, z7  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11;
  output z0, z1, z2, z3, z4, z5, z6, z7;
  assign z0 = ~x02 & ((x04 & ((~x08 & (x00 ? ~x07 : (~x01 & ~x03 & x06 & x10 & ((x11 & ((x05 & (x07 ^ x09)) | (x07 & x09))) | (~x05 & x07 & ~x09))))) | (~x00 & ~x01 & ~x03 & ~x06 & x10 & (x05 ? x11 : (~x09 | (x09 & x11)))))) | (~x00 & ~x01 & ~x03 & ~x04));
  assign z1 = ~x02 & x04 & (x00 ? (x07 & x08) : (~x01 & ~x03 & ~x10 & ((x11 & (x06 ? (~x08 & ((x05 & (x07 ^ x09)) | (x07 & x09))) : (x05 | (~x05 & x09)))) | (~x05 & ~x09 & (~x06 | (x06 & x07 & ~x08))))));
  assign z2 = ~x02 & x04 & (x00 ? (x07 & ~x08) : (~x01 & ~x03 & ((x09 & ((~x05 & (x06 ? (~x07 & ~x08) : ~x11)) | (x06 & ~x08 & ~x11 & (x07 | (x05 & ~x07))))) | (x05 & (x06 ? (~x08 & ~x09 & (~x07 | (x07 & ~x11))) : ~x11)))));
  assign z3 = x00 ? (~x04 & ~x08 & (~x07 | (x02 & x07))) : (~x01 & ~x02 & ~x03 & x04 & x06 & ((x08 & ((x05 & (~x07 | (x07 & x09))) | (x07 & ~x09) | (~x05 & x09))) | (~x05 & ~x07 & ~x09)));
  assign z4 = (x00 & ~x04 & x08 & (~x07 | (x02 & x07))) | (~x00 & ~x01 & ~x02 & x03);
  assign z5 = (~x00 & ~x01 & x02) | (x00 & ~x02 & ~x04 & x07 & ~x08);
  assign z6 = (~x00 & x01) | (x00 & ~x02 & ~x04 & x07 & x08);
  assign z7 = x00 & x04 & ((x02 & (~x08 | (x07 & x08))) | (~x07 & x08));
endmodule