module pla__in1 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16;
  assign z00 = (~x13 & (x10 ? (x11 ? ((~x00 & ((~x06 & ((~x14 & ((~x08 & ((x04 & ~x05 & x12 & (x09 | (x07 & ~x09))) | (x07 & ~x12 & ~x15))) | (x05 & ~x12))) | (~x12 & ((~x07 & ~x15 & (x08 | x09)) | (x05 & x08))))) | (x05 & ~x12 & (~x15 | (x08 & ~x14))))) | (x05 & x06 & x07 & ~x12 & (~x15 | (x08 & ~x14)))) : (x12 ? ((x00 & (x15 ? ~x01 : ~x14)) | x14 | (~x00 & ~x14 & x15)) : ((x04 & ~x05 & ~x06 & x07 & ~x14 & (x08 | (~x08 & x09)) & (~x00 | ~x15)) | (~x00 & x14)))) : (x04 ? (x11 ? ((x05 & ((~x00 & ((x01 & ((x06 & ~x14 & x15) | (~x12 & ~x15 & ~x06 & x08))) | (~x14 & ((x06 & x15 & (x07 | (~x01 & ~x07 & x12))) | (~x12 & ~x15 & (~x06 | (~x07 & x08))))) | (~x12 & x14 & x15 & (~x06 | (~x07 & x08))))) | (x06 & x07 & x08 & ~x12 & (x14 ^ ~x15)))) | (~x07 & x08 & ~x05 & ~x06 & ~x14 & ~x15 & x09 & x12)) : (x12 & (~x15 | (x15 & (x14 | (~x06 & ~x14)))))) : (~x11 & (x12 | (~x05 & ~x14)))))) | (x13 & ((x12 & ((x04 & ((~x00 & x05 & ~x10 & x11 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14))) | (~x14 & x15 & x10 & ~x11))) | (x10 & ~x11 & ((x14 & ~x15) | (~x04 & ~x14 & x15 & (x07 | (~x07 & ((~x06 & ~x08 & x09) | (x08 & ~x09))))))) | (~x05 & ~x10 & x11 & ~x14))) | (~x12 & ((x04 & ((~x05 & ~x06 & ~x07 & x11 & x15 & ((~x08 & x09 & x14) | (x08 & ~x09 & ~x10 & ~x14))) | (~x10 & ~x11))) | (x10 & ~x11 & (~x14 | (x14 & ((x07 & ~x08 & x09) | (x08 & ~x15))))))) | (~x14 & ~x15 & x10 & ~x11))) | (~x04 & ~x10 & ~x11 & ~x12 & ~x15);
  assign z01 = (~x13 & (x11 ? ((~x00 & ((x05 & (x10 ? (~x12 & (~x15 | (x08 & ~x14) | (~x06 & (x08 | ~x14)))) : ((~x14 & ((x06 & x15 & (((~x04 | (x04 & x09)) & (x01 | x07)) | (x12 & (~x04 | (~x01 & x04 & ~x07 & x09))))) | (~x04 & ~x12 & ~x15 & (~x06 | x08)))) | (~x04 & ~x12 & x14 & x15 & (~x06 | x08))))) | (~x06 & x10 & ((~x12 & ~x15 & (x07 ? (~x08 & ~x14) : (x08 | x09))) | (~x05 & ~x08 & x12 & ~x14 & (x09 | (x07 & (~x04 | (x04 & ~x09))))))))) | (~x10 & ((~x07 & x08 & ~x05 & ~x06 & ~x14 & ~x15 & x09 & x12) | (~x12 & ((~x04 & ((x14 & ~x15) | (x05 & x06 & x07 & x08 & (x14 ^ ~x15)))) | (x14 & ~x15 & (x06 | ~x08 | ~x01 | ~x05)))))) | (x05 & x06 & x07 & x10 & ~x12 & (~x15 | (x08 & ~x14)))) : (x10 ? (x12 ? (x00 ? (x15 ? ~x01 : ~x14) : (~x14 & x15)) : ((~x00 & x14) | (~x05 & ~x06 & x07 & ~x14 & (~x00 | ~x15) & (x08 | (x09 & (~x04 | (x04 & ~x08))))))) : ((~x01 & ~x12 & x14 & (x00 | x15)) | x12 | (~x04 & ~x05 & ~x14))))) | (x13 & ((~x14 & ((x12 & (x10 ? (~x11 & x15 & (x04 | (~x04 & (x07 | (~x07 & ((~x06 & ~x08 & x09) | (x08 & ~x09))))))) : (x11 & (~x05 | (~x00 & ~x02 & x05 & x06 & (~x04 | (x04 & x09)) & (x01 | x07)))))) | (x10 & ~x11 & (~x12 | ~x15)) | (~x07 & x08 & ~x05 & ~x06 & ~x09 & ~x10 & x11 & ~x12 & x15))) | (x05 & ~x10 & ((~x11 & ~x12 & x15) | (~x00 & x01 & ~x04 & ~x06 & x08 & x11 & x12 & x14 & ~x15))) | (x14 & ((~x12 & ((~x08 & x09 & ((x07 & x10 & ~x11) | (~x05 & ~x06 & ~x07 & x11 & x15))) | (x08 & x10 & ~x11 & ~x15))) | (x10 & ~x11 & x12))))) | (~x10 & ~x11 & ~x12 & (x04 | (x05 & ~x14 & x15) | (~x04 & ~x15)));
  assign z02 = (~x13 & (x11 ? ((~x10 & ((~x07 & x08 & ~x05 & ~x06 & ~x14 & ~x15 & x09 & x12) | (~x12 & ((~x04 & ((x14 & ~x15) | (x05 & x06 & x07 & x08 & (x14 ^ ~x15)))) | (x14 & ~x15 & (x06 | ~x08 | ~x01 | ~x05)))))) | (x05 & x06 & x07 & x10 & ~x12 & (~x15 | (x08 & ~x14))) | (~x00 & ((x05 & (x10 ? (~x12 & (~x15 | (x08 & ~x14) | (~x06 & (x08 | ~x14)))) : ((x01 & ((x06 & ~x14 & x15) | (x04 & ~x06 & x08 & ~x12 & ~x15))) | (~x04 & ((~x12 & (x14 ^ ~x15) & (~x06 | x08)) | (~x14 & x15 & x06 & x12))) | (x06 & ~x14 & x15 & (x07 | (~x07 & x12 & ~x01 & x04)))))) | (~x06 & x10 & ((~x08 & ~x14 & ((x07 & ~x12 & ~x15) | (~x05 & x12 & (x07 | (~x04 & x09))))) | (~x07 & ~x12 & ~x15 & (x08 | x09))))))) : ((x00 & ((~x01 & ~x10 & ~x12 & x14) | (~x14 & ~x15 & x10 & x12))) | (x10 & ((~x12 & ((~x00 & x14) | (~x05 & ~x06 & x07 & ~x14 & (~x00 | ~x15) & (x08 | (x09 & (~x04 | (x04 & ~x08))))))) | (~x14 & x15 & ~x00 & x12))) | (~x10 & (x12 | (~x04 & ~x05 & ~x14) | (x14 & x15 & ~x01 & ~x12)))))) | (x13 & ((x12 & (x10 ? (~x11 & ~x14 & x15 & (x04 | (~x04 & (x07 | (~x07 & ((~x06 & ~x08 & x09) | (x08 & ~x09))))))) : (x11 & ((~x05 & ~x14) | (~x00 & x05 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14))))))) | (~x14 & ~x15 & x10 & ~x11) | (~x12 & ((x15 & (x05 ? (~x10 & ~x11) : (~x06 & ~x07 & x11 & ((x08 & ~x09 & ~x10 & ~x14) | (x09 & x14 & ~x04 & ~x08))))) | (x10 & ~x11 & x14 & ((x07 & ~x08 & x09) | (x08 & ~x15))))))) | (~x11 & (x10 ? (x12 & x14) : (~x12 & (x04 | (x05 & ~x14 & x15) | (~x04 & ~x15)))));
  assign z03 = x11 ? ((~x10 & ((x05 & ((~x00 & ((~x14 & ((x06 & (((x01 | x07) & ((~x02 & x12 & x13) | (~x13 & x15))) | (~x13 & x15 & ~x04 & x12))) | (~x12 & ~x13 & ~x15 & (~x06 | (x08 & (~x04 | (x04 & ~x07))))))) | (~x06 & ((x01 & x08 & ~x15 & ((x04 & ~x12 & ~x13) | (x12 & x13 & x14))) | (~x04 & ~x12 & ~x13 & x14 & x15))) | (~x13 & x14 & x15 & ~x04 & x08 & ~x12))) | (x06 & x07 & x08 & ~x12 & ~x13 & ((~x14 & ~x15) | (~x04 & x14 & x15))))) | (~x05 & ((~x14 & ((x12 & x13) | (~x06 & ~x07 & x08 & ((~x09 & ~x12 & x13 & x15) | (x09 & x12 & ~x13 & ~x15))))) | (x14 & ~x15 & ~x12 & ~x13))) | (~x12 & ~x13 & x14 & ~x15 & (x06 | ~x08 | ~x01 | ~x04)))) | (~x06 & ((~x08 & ((~x05 & ((~x00 & x10 & x12 & ~x13 & ~x14 & (x07 | (~x04 & x09))) | (~x04 & ~x07 & x09 & x14 & x15 & ~x12 & x13))) | (~x00 & x07 & x10 & ~x14 & ~x15 & ~x12 & ~x13))) | (~x00 & x10 & ~x12 & ~x13 & ((~x07 & ~x15 & (x08 | x09)) | (x05 & (x08 | ~x14)))))) | (x05 & x10 & ~x12 & ~x13 & (~x15 | (x08 & ~x14)) & (~x00 | (x06 & x07)))) : ((~x12 & (x10 ? ((x07 & ((~x05 & ~x06 & ~x13 & ~x14 & (~x00 | ~x15) & (x08 | (x09 & (~x04 | (x04 & ~x08))))) | (~x08 & x09 & x13 & x14))) | (x13 & (~x14 | (x08 & x14 & ~x15))) | (~x00 & ~x13 & x14)) : ((x15 & ((~x13 & x14) ? ~x01 : x05)) | x04 | (~x01 & ~x13 & x14 & (x00 | (~x00 & ~x04 & ~x15)))))) | (x12 & (x10 ? (x13 ? (x15 & (x14 | (~x14 & (x04 | (~x04 & (x07 | (~x07 & ((~x06 & ~x08 & x09) | (x08 & ~x09))))))))) : ((x00 & (x15 ? ~x01 : ~x14)) | x14 | (~x00 & ~x14 & x15))) : (~x13 & (x04 | (~x14 & x15 & ~x01 & x06))))) | (~x14 & ~x15 & x10 & x13));
  assign z04 = x11 ? ((~x00 & ((x05 & (x10 ? (~x12 & ~x13 & (~x15 | (x08 & ~x14) | (~x06 & (x08 | ~x14)))) : ((~x14 & ((x06 & (((x01 | x07) & ((~x02 & x12 & x13) | (~x13 & x15))) | (~x13 & x15 & ~x04 & x12))) | (~x04 & ~x12 & ~x13 & ~x15 & (~x06 | x08)))) | (~x04 & x14 & ((~x06 & ((~x12 & ~x13 & x15) | (x01 & x08 & x12 & x13 & ~x15))) | (~x13 & x15 & x08 & ~x12)))))) | (~x06 & x10 & ~x13 & ((~x12 & ~x15 & (x07 ? (~x08 & ~x14) : (x08 | x09))) | (~x05 & ~x08 & x12 & ~x14 & (x09 | (x07 & (~x04 | (x04 & ~x09))))))))) | (~x12 & ((~x05 & ((~x06 & ~x07 & x13 & x15 & ((~x08 & x09 & x14) | (x08 & ~x09 & ~x10 & ~x14))) | (x14 & ~x15 & ~x10 & ~x13))) | (~x13 & ((x06 & ((x05 & x07 & ((x10 & (~x15 | (x08 & ~x14))) | (x08 & ~x10 & (x14 ^ ~x15)))) | (~x10 & x14 & ~x15))) | (~x10 & x14 & ~x15 & (~x01 | ~x04 | ~x08)))))) | (~x05 & ~x10 & x12 & ~x14 & (x13 | (~x06 & ~x07 & x08 & x09 & ~x13 & ~x15)))) : ((~x12 & ((~x13 & ((x14 & ((~x01 & ~x10 & (x00 | x15)) | (~x00 & x10))) | (~x05 & ~x06 & x07 & x10 & ~x14 & (~x00 | ~x15) & (x08 | (x09 & (~x04 | (x04 & ~x08))))))) | (~x10 & ((x05 & x15 & (x13 | ~x14)) | x04 | (~x04 & ~x15))) | (x10 & x13 & (~x14 | (x14 & ((x07 & ~x08 & x09) | (x08 & ~x15))))))) | (x12 & (x10 ? (x13 ? (x14 | (~x14 & x15 & (x04 | (~x04 & (x07 | (~x07 & ((~x06 & ~x08 & x09) | (x08 & ~x09)))))))) : (x00 ? (x15 ? ~x01 : ~x14) : (~x14 & x15))) : ~x13)) | (~x04 & ~x05 & ~x10 & ~x13 & ~x14));
  assign z05 = ~x11 & ((~x12 & ((x10 & x13 & ~x14) | (~x04 & ~x10 & ~x15))) | (~x13 & ((~x04 & ~x10 & (x12 | (~x05 & ~x14))) | (x00 & ~x01 & x10 & x12 & x15))) | (x10 & ((x12 & x14) | (x13 & ~x14 & ~x15))));
  assign z06 = x10 ? ((~x13 & (x11 ? (~x12 & ((x05 & (((~x15 | (x08 & ~x14)) & (~x00 | (x06 & x07))) | (~x00 & ~x06 & (x08 | ~x14)))) | (~x00 & ~x06 & ~x15 & (x07 ? (~x08 & ~x14) : (x08 | x09))))) : (x12 & (x00 ? (x15 ? ~x01 : ~x14) : (~x14 & x15))))) | (~x11 & ((x12 & x14) | (x13 & ((~x14 & ~x15) | (~x12 & (~x14 | (x14 & ((x07 & ~x08 & x09) | (x08 & ~x15)))))))))) : (~x11 & ((~x12 & ((~x04 & ~x15) | (x14 & x15 & x04 & x13))) | (~x13 & (x04 ? (x12 & (~x15 | (x15 & (x14 | (~x06 & ~x14))))) : (x12 | (~x05 & ~x14))))));
  assign z07 = (~x13 & (x11 ? ((~x10 & ((x05 & ((x06 & x07 & x08 & ~x12 & (x14 ^ ~x15)) | (~x00 & ((x01 & ((x06 & ~x14 & x15) | (x04 & ~x06 & x08 & ~x12 & ~x15))) | (~x12 & (x14 ^ ~x15) & (~x06 | (x08 & (~x04 | (x04 & ~x07))))) | (x06 & ~x14 & x15 & (x07 | (x12 & (~x04 | (~x01 & x04 & ~x07))))))))) | (~x15 & ((~x05 & ((~x12 & x14) | (~x06 & ~x07 & x08 & x09 & x12 & ~x14))) | (~x12 & x14 & (x06 | ~x08 | ~x01 | ~x04)))))) | (~x00 & ~x05 & ~x06 & ~x08 & x10 & x12 & ~x14 & (x09 | (x07 & (~x04 | (x04 & ~x09)))))) : ((~x01 & ((x00 & (x10 ? (x12 & x15) : (~x12 & x14))) | (~x10 & x15 & ((~x12 & x14) | (x06 & x12 & ~x14))))) | (~x12 & (x10 ? ((~x00 & x14) | (~x05 & ~x06 & x07 & ~x14 & (~x00 | ~x15) & (x08 | (x09 & (~x04 | (x04 & ~x08)))))) : x04)) | (~x10 & ((~x04 & (x12 | (~x05 & ~x14))) | (x04 & x06 & x12 & ~x14 & x15)))))) | (x13 & ((~x10 & (x11 ? ((x12 & ((~x05 & ~x14) | (~x00 & x05 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14))))) | (~x07 & x08 & ~x05 & ~x06 & ~x14 & x15 & ~x09 & ~x12)) : (~x12 & ((x04 & (~x15 | (~x14 & x15))) | (x05 & x15))))) | (x15 & ((~x07 & ((~x04 & x10 & ~x11 & x12 & ~x14 & ((~x06 & ~x08 & x09) | (x08 & ~x09))) | (~x05 & ~x06 & ~x08 & ~x12 & x14 & x09 & x11))) | (x10 & ~x11 & x12 & ~x14 & (x04 | (~x04 & x07))))) | (x10 & ~x11 & ~x14 & (~x12 | ~x15)))) | (~x11 & (x10 ? (x12 & x14) : (~x12 & ((x05 & ~x14 & x15) | (~x04 & ~x15)))));
  assign z08 = (~x13 & ((x12 & (x10 ? (x00 ? (~x11 & (x15 ? ~x01 : ~x14)) : (x04 & ~x05 & ~x06 & ~x08 & x11 & ~x14 & (x09 | (x07 & ~x09)))) : (x04 ? (~x07 & x11 & ~x14 & ((~x00 & ~x01 & x05 & x06 & x15) | (~x05 & ~x06 & x08 & x09 & ~x15))) : ~x11))) | (x04 & (x05 ? (~x10 & x11 & ((x06 & x07 & x08 & ~x12 & (x14 ^ ~x15)) | (~x00 & ((x01 & ((x06 & ~x14 & x15) | (~x12 & ~x15 & ~x06 & x08))) | (~x12 & (~x06 | (~x07 & x08)) & (x14 ^ ~x15)) | (~x14 & x15 & x06 & x07))))) : (~x06 & x07 & ~x08 & x09 & x10 & ~x11 & ~x12 & ~x14 & (~x00 | ~x15)))) | (~x04 & ~x05 & ~x10 & ~x11 & ~x14))) | (x13 & ((x04 & ((~x10 & (x11 ? ((~x07 & x08 & ~x05 & ~x06 & ~x14 & x15 & ~x09 & ~x12) | (~x00 & x05 & x12 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14)))) : (~x12 & (~x15 | (~x14 & x15))))) | (~x05 & ~x06 & ~x07 & ~x08 & x09 & x11 & ~x12 & x14 & x15))) | (x10 & ~x11 & ((~x14 & ~x15) | (~x12 & (~x14 | (x14 & ((x07 & ~x08 & x09) | (x08 & ~x15))))))) | (~x05 & ~x10 & x11 & x12 & ~x14))) | (~x11 & ((x10 & x12 & x14) | (~x12 & ~x15 & ~x04 & ~x10)));
  assign z09 = (~x13 & ((x04 & ((~x06 & ~x14 & ((~x05 & ((x10 & ((~x00 & ((~x07 & ~x08 & x09 & x11 & x12) | (x07 & x08 & ~x11 & ~x12))) | (~x11 & ~x12 & ~x15 & x07 & x08))) | (~x07 & x08 & x09 & ~x10 & x11 & x12 & ~x15))) | (~x10 & ~x11 & x12 & x15))) | (~x10 & ~x11 & x12 & x14))) | (~x11 & ((~x04 & ~x10 & (x12 | (~x05 & ~x14))) | (x00 & ~x01 & x10 & x12 & x15))))) | (~x04 & ~x10 & ~x11 & ~x12 & ~x15) | (x10 & ((x13 & ((~x11 & ~x14 & (~x12 | ~x15)) | (x09 & x11 & ~x12 & x14 & x15 & x04 & ~x05 & ~x06 & ~x07 & ~x08))) | (~x11 & x12 & x14)));
  assign z10 = x10 ? ((~x11 & ((x12 & ((x00 & ~x13 & (x15 ? ~x01 : ~x14)) | x14 | (x13 & ~x14 & x15 & (x04 | (~x04 & x07 & ~x08))))) | (x13 & ~x14 & ~x15) | (~x12 & ((~x00 & ~x13 & x14) | (x13 & ~x14))))) | (~x00 & x04 & ~x05 & ~x06 & x07 & ~x08 & ~x09 & x11 & x12 & ~x13 & ~x14)) : ((~x12 & ((~x13 & ((x14 & ((x15 & ((x04 & x05 & x11 & ((~x00 & (~x06 | (~x07 & x08))) | (x06 & x07 & x08))) | (~x01 & ~x11))) | (x00 & ~x01 & ~x11))) | (x04 & x05 & x11 & ~x15 & ((~x00 & ((~x06 & (~x14 | (x01 & x08))) | (~x07 & x08 & ~x14))) | (x08 & ~x14 & x06 & x07))))) | (~x11 & ((x05 & x15 & (x13 | ~x14)) | x04 | (~x04 & ~x15))) | (x04 & ~x05 & ~x06 & ~x07 & x11 & x13 & x15 & (x08 ? (~x09 & ~x14) : (x09 & x14))))) | (~x00 & x04 & x05 & x11 & ((x06 & ~x14 & (x01 | x07) & ((~x02 & x12 & x13) | (~x13 & x15))) | (x01 & ~x06 & x08 & x14 & ~x15 & x12 & x13))) | (~x04 & ~x11 & ~x13 & (x12 | (~x05 & ~x14))));
  assign z11 = x11 ? ((~x06 & ((~x00 & x12 & ((x04 & ~x05 & ~x08 & ~x13 & ~x14 & x09 & x10) | (x05 & x08 & x01 & ~x04 & x14 & ~x15 & ~x10 & x13))) | (x04 & ~x05 & ~x07 & ~x08 & x09 & x10 & ~x12 & x13 & x14 & x15))) | (~x10 & ((~x12 & ~x13 & x14 & ~x15 & (x06 | ~x08 | ~x01 | ~x04)) | (~x05 & ((x14 & ~x15 & ~x12 & ~x13) | (x12 & x13 & ~x14)))))) : (x10 ? ((~x13 & ((~x12 & ((x04 & ~x05 & ~x06 & x07 & ~x14 & (x08 | (~x08 & x09)) & (~x00 | ~x15)) | (~x00 & x14))) | (x00 & x12 & (x15 ? ~x01 : ~x14)))) | (x12 & x14) | (x13 & ((x07 & ((~x08 & x09 & ~x12 & x14) | (x12 & ~x14 & x15 & ~x04 & x08))) | (~x14 & (~x12 | ~x15 | (~x04 & ~x07 & x12 & x15 & ((~x06 & ~x08 & x09) | (x08 & ~x09))))) | (x14 & ~x15 & x08 & ~x12)))) : ((~x13 & ((~x04 & (x12 | (~x05 & ~x14))) | (x06 & x12 & ~x14 & x15 & (~x01 | x04)))) | (~x12 & (x04 ? (x13 & (~x15 | (~x14 & x15))) : ~x15))));
  assign z12 = x11 ? (x13 ? ((~x10 & ((x12 & ((~x00 & ~x04 & x05 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14))) | (~x05 & ~x14 & ~x15))) | (~x05 & ~x06 & ~x07 & ~x12 & x15 & ((x08 & ~x09 & ~x14) | (x09 & x14 & x04 & ~x08))))) | (~x04 & ~x05 & ~x06 & ~x07 & ~x08 & x09 & ~x12 & x14 & x15)) : ((~x00 & ((x05 & (x10 ? (~x12 & (~x15 | (x08 & ~x14) | (~x06 & (x08 | ~x14)))) : ((x01 & ((x04 & ~x06 & x08 & ~x12 & ~x15) | (~x14 & x15 & ~x04 & x06))) | (~x12 & (x14 ^ ~x15) & (~x06 | (x08 & (~x04 | (x04 & ~x07))))) | (x06 & ~x14 & x15 & ((~x07 & x12 & ~x01 & x04) | (~x04 & (x07 | x12))))))) | (~x06 & x10 & ((~x07 & ~x12 & ~x15 & (x08 | x09)) | (~x08 & ~x14 & ((x07 & ~x12 & ~x15) | (~x05 & x12 & (x04 ? (x07 & x09) : (x07 | x09))))))))) | (x05 & x06 & x07 & x10 & ~x12 & (~x15 | (x08 & ~x14))) | (~x10 & ((~x15 & ((~x04 & ((~x12 & x14) | (~x05 & ~x06 & ~x07 & x12 & ~x14 & x08 & x09))) | (~x12 & ((x06 & (x14 | (x08 & ~x14 & x05 & x07))) | (x14 & (~x01 | ~x05 | ~x08)))))) | (x05 & x06 & x07 & x14 & x15 & x08 & ~x12))))) : ((~x13 & ((x12 & ((x15 & ((~x01 & ((x00 & x10) | (x06 & ~x10 & ~x14))) | (~x00 & x10 & ~x14))) | (~x10 & (~x04 | (x04 & ~x14))))) | (~x05 & ~x14 & ((~x04 & ~x10) | (~x06 & x07 & x10 & ~x12 & (~x00 | ~x15) & (x08 | (x09 & (~x04 | (x04 & ~x08))))))))) | (~x12 & (x10 ? (x13 & ~x14) : (x04 ? (x13 & x15) : ~x15))) | (x10 & ((x13 & ~x14 & ~x15) | (x12 & (x14 | (~x04 & x13 & ~x14 & x15 & ((x08 & ~x09) | (~x08 & x09 & ~x06 & ~x07))))))));
  assign z13 = (~x13 & (x11 ? ((~x00 & ((~x14 & (x05 ? (~x10 & ((~x04 & ~x12 & ~x15 & (~x06 | x08)) | (x06 & x15 & ((~x04 & x12) | ((x01 | x07) & (~x04 | (x04 & ~x09))))))) : (~x06 & ~x08 & x10 & x12 & (x04 ? (x07 & x09) : (x07 | x09))))) | (~x04 & x05 & ~x10 & ~x12 & x14 & x15 & (~x06 | x08)))) | (x08 & ~x10 & ((~x04 & x05 & x06 & x07 & ~x12 & (x14 ^ ~x15)) | (~x14 & ~x15 & x09 & x12 & ~x05 & ~x06 & ~x07)))) : (x10 ? ((x00 & x12 & (x15 ? ~x01 : ~x14)) | (~x05 & ~x06 & x07 & ~x12 & ~x14 & (~x00 | ~x15) & (x04 ? (~x08 & x09) : (x08 | x09)))) : ((~x04 & ~x05 & ~x14) | (x12 & (~x04 | (x04 & ((x14 & ~x15) | (~x06 & ~x14 & x15))))))))) | (~x11 & ((x10 & x12 & x14) | (~x12 & ~x15 & ~x04 & ~x10))) | (x13 & (x11 ? ((~x04 & ~x05 & ~x06 & ~x07 & ~x08 & x09 & ~x12 & x14 & x15) | (~x10 & ((~x14 & ((x12 & ((~x00 & ~x02 & x05 & x06 & (x01 | x07) & (~x04 | (x04 & ~x09))) | (~x05 & x15))) | (~x04 & ~x05 & ~x06 & ~x07 & x08 & ~x09 & ~x12 & x15))) | (~x00 & x01 & x04 & x05 & ~x06 & x08 & ~x09 & x12 & x14 & ~x15)))) : ((~x12 & ((x10 & ~x14) | (x04 & ~x10 & ~x15))) | (x10 & ~x14 & (~x15 | (~x04 & x07 & x08 & ~x09 & x12 & x15))))));
  assign z14 = (~x10 & (x11 ? (x13 ? ((~x05 & ~x06 & ~x07 & ~x12 & x15 & ((x08 & ~x09 & ~x14) | (x09 & x14 & x04 & ~x08))) | (x12 & ((~x00 & x05 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14)) & (~x04 | (x04 & x09))) | (~x05 & ~x14 & x15)))) : ((~x01 & ((~x00 & x04 & x05 & x06 & x12 & ~x14 & x15 & ~x07 & ~x09) | (~x12 & x14 & ~x15))) | (~x15 & ((~x05 & ~x06 & ~x07 & x12 & ~x14 & x08 & x09) | (~x12 & ((x05 & ((x08 & ~x14 & x06 & x07) | (~x00 & ((~x06 & ~x14) | (x08 & (x04 ? ((x01 & ~x06) | (~x07 & ~x14)) : ~x14)))))) | (x14 & (x06 | ~x08 | ~x04 | ~x05)))))) | (x05 & x15 & ((~x00 & ((x06 & ~x14 & (((~x04 | (x04 & x09)) & (x01 | x07)) | (~x04 & x12))) | (~x12 & x14 & (~x06 | (x08 & (~x04 | (x04 & ~x07))))))) | (x06 & x07 & x08 & ~x12 & x14))))) : ((x04 & (x12 ? (~x13 & (x14 | (~x14 & x15))) : (x13 & (~x14 | (x14 & x15))))) | (~x13 & ((~x04 & (x12 | (~x05 & ~x14))) | (~x01 & x06 & x12 & ~x14 & x15))) | (~x04 & ~x12 & ~x15)))) | (x13 & ((x10 & ~x11 & ((~x14 & ~x15) | (~x12 & (~x14 | (x14 & ((x07 & ~x08 & x09) | (x08 & ~x15))))))) | (x15 & ((~x04 & ((~x06 & ~x07 & ~x08 & x09 & ((~x12 & x14 & ~x05 & x11) | (x10 & ~x11 & x12 & ~x14))) | (x08 & ~x09 & x10 & ~x11 & x12 & ~x14))) | (~x11 & x12 & ~x14 & x04 & x10))))) | (x10 & ((~x11 & ((x12 & x14) | (~x13 & ((~x12 & ((~x00 & (x14 | (x04 & ~x05 & ~x06 & x07 & x09 & ~x14))) | (x04 & ~x05 & ~x06 & ~x14 & ~x15 & x07 & x09))) | (x12 & x15 & x00 & ~x01))))) | (~x00 & ~x05 & ~x06 & ~x08 & x11 & x12 & ~x13 & ~x14 & (x09 | (x07 & (~x04 | (x04 & ~x09 & ~x15)))))));
  assign z15 = (~x13 & (x11 ? ((~x00 & ((x05 & ((x10 & ~x12 & (~x15 | (x08 & ~x14) | (~x06 & (x08 | ~x14)))) | (x04 & ~x10 & ((x01 & ((~x12 & ~x15 & ~x06 & x08) | (~x14 & x15 & x06 & x09))) | (~x12 & x14 & x15 & (~x06 | (~x07 & x08))) | (~x14 & ((~x12 & ~x15 & (~x06 | (~x07 & x08))) | (x06 & x09 & x15 & (x07 | (~x01 & ~x07 & x12))))))))) | (~x06 & x10 & ((~x07 & ~x12 & ~x15 & (x08 | x09)) | (~x08 & ~x14 & ((x07 & ~x12 & ~x15) | (~x05 & x09 & x12 & (~x04 | (x04 & x07))))))))) | (x05 & x06 & x07 & ~x12 & ((x08 & ((x10 & ~x14) | (x04 & ~x10 & (x14 ^ ~x15)))) | (x10 & ~x15)))) : ((~x01 & ((x00 & (x10 ? (x12 & x15) : (~x12 & x14))) | (x14 & x15 & ~x10 & ~x12))) | (~x10 & (x04 ? (~x12 | (x12 & ((x14 & ~x15) | (~x06 & ~x14 & x15)))) : (x12 | (~x05 & ~x14)))) | (x10 & ~x12 & ((~x00 & x14) | (x04 & ~x05 & ~x06 & x07 & ~x14 & (~x00 | ~x15) & (x08 ^ x09))))))) | (~x11 & (x10 ? (x12 & x14) : (~x12 & ((x05 & ~x14 & x15) | (~x04 & ~x15))))) | (x13 & ((x12 & ((x04 & ((~x14 & x15 & x10 & ~x11) | (~x00 & x05 & x09 & ~x10 & x11 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14))))) | (~x14 & x15 & ((~x04 & x10 & ~x11 & (x07 ? (~x08 | (x08 & x09)) : (x08 & ~x09))) | (~x05 & ~x10 & x11))))) | (~x14 & ~x15 & x10 & ~x11) | (~x12 & (x10 ? (~x11 & ~x14) : (x15 & ((x04 & x14 & (~x11 | (~x05 & ~x06 & ~x07 & ~x08 & x09 & x11))) | (x05 & ~x11)))))));
  assign z16 = (~x13 & (x10 ? (x11 ? ((x05 & x06 & x07 & ~x12 & (~x15 | (x08 & ~x14))) | (~x00 & ((x05 & ~x12 & (~x15 | (x08 & ~x14))) | (~x06 & ((~x12 & ((~x07 & ~x15 & (x08 | x09)) | (x05 & x08))) | (~x14 & ((x05 & ~x12) | (~x08 & ((x07 & ~x12 & ~x15) | (~x05 & x12 & (x04 ? (x07 ? (~x09 & x15) : x09) : (x07 | x09)))))))))))) : (x12 ? (x00 ? (x15 ? ~x01 : ~x14) : (~x14 & x15)) : ((~x00 & x14) | (~x05 & ~x06 & x07 & ~x14 & (~x00 | ~x15) & (x04 ? (x08 & ~x09) : (x08 | x09)))))) : ((~x01 & ((x12 & ~x14 & x15 & x06 & ~x11) | (x14 & ~x15 & x11 & ~x12))) | (~x14 & ((x12 & ((x04 & ~x11 & (~x15 | (x06 & x15))) | (x11 & ((x05 & x06 & x15 & ~x00 & ~x04) | (x08 & x09 & ~x15 & ~x05 & ~x06 & ~x07))))) | (~x04 & (x05 ? (x11 & ((x06 & ((~x00 & x15 & (x01 | x07)) | (~x12 & ~x15 & x07 & x08))) | (~x00 & ~x12 & ~x15 & (~x06 | x08)))) : ~x11)))) | (x14 & ((x11 & ~x12 & ((~x04 & (~x15 | (x05 & x15 & ((x06 & x07 & x08) | (~x00 & (~x06 | x08)))))) | (~x15 & (~x05 | x06 | ~x08)))) | (x12 & x15 & x04 & ~x11))) | (~x04 & ~x11 & x12)))) | (~x11 & ((x10 & x12 & x14) | (~x12 & ~x15 & ~x04 & ~x10))) | (x13 & ((~x10 & ((x11 & ((~x07 & x08 & ~x05 & ~x06 & ~x14 & x15 & ~x09 & ~x12) | (x12 & ((~x00 & ~x04 & x05 & ((x01 & ((~x02 & x06 & ~x14) | (~x06 & x08 & x14 & ~x15))) | (~x02 & x06 & x07 & ~x14))) | (~x05 & ~x14 & ~x15))))) | (x04 & ~x11 & ~x12 & (x14 | (~x14 & x15))))) | (~x12 & ((x10 & ~x11 & ~x14) | (x14 & ((x08 & x10 & ~x11 & ~x15) | (~x08 & x09 & ((x07 & x10 & ~x11) | (~x05 & ~x06 & ~x07 & x11 & x15 & (~x04 | (x04 & x10))))))))) | (x10 & ~x11 & ~x14 & (~x15 | (~x04 & ~x07 & x12 & x15 & ((~x06 & ~x08 & x09) | (x08 & ~x09)))))));
endmodule