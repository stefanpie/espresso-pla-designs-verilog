module pla__sao2 ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,
    z0, z1, z2, z3  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output z0, z1, z2, z3;
  assign z0 = ~x5 & ~x9 & ((x7 & ((~x4 & ((x1 & x3 & x8 & (x6 ? ~x2 : x0)) | (~x1 & ~x2 & ~x3 & ~x6 & ~x8))) | (x0 & x2 & ((~x1 & x4 & (x3 ? ~x8 : x6)) | (~x6 & ~x8 & x1 & x3))))) | (~x0 & x3 & ((x1 & x4 & x6 & x8 & (~x2 | ~x7)) | (~x2 & ~x4 & ~x6 & ~x8 & (~x1 | ~x7)))));
  assign z1 = ~x5 & ~x9 & (((~x1 ^ x8) & ((x0 & x7 & ((x2 & x4 & (x3 ^ x6)) | (~x2 & x3 & ~x4 & ~x6))) | (~x0 & ~x2 & x3 & ~x4 & ~x6 & ~x7))) | ((~x0 ^ x2) & ((x1 & x3 & ((~x4 & x7 & (x6 ^ ~x8)) | (x4 & x6 & ~x7 & x8))) | (~x1 & ~x3 & ~x4 & ~x6 & x7 & ~x8))) | (x3 & x4 & x6 & x7 & ((x0 & (x1 ? (x2 ^ x8) : (x2 & x8))) | (x2 & x8 & ~x0 & x1))));
  assign z2 = ~x9 & ((~x5 & (((~x0 | ~x7) & ((x2 & ~x4) | (~x1 & x8) | (x6 & ~x8))) | (~x6 & ((~x1 & x8) | (x4 & (~x2 | ~x7)))) | ((~x2 | ~x4) & ((~x1 & x8) | (x6 & ~x8) | (x1 & ~x3))) | (x1 & ~x3 & (~x0 | ~x8)) | (x0 & ~x2 & ~x7))) | (~x3 & (~x7 | (x1 & ~x6))) | x5 | (~x0 & x4 & ~x6));
  assign z3 = ~x5 & ~x9 & ((x0 & ((~x2 & ~x7) | (~x1 & x2 & ~x3 & ~x4 & ~x6 & x7 & ~x8))) | ((~x0 | ~x7) & ((~x1 & x8) | (x6 & ~x8) | (x2 & ~x4) | (x1 & ~x3))) | ((~x2 | ~x4) & ((~x1 & x8) | (x6 & ~x8) | (x1 & ~x3))) | (~x7 & (x4 ? ~x6 : x3)) | (~x6 & ((~x1 & (x8 | (~x2 & ~x3 & ~x4 & x7 & ~x8))) | (x4 & (~x2 | ~x3)) | (~x0 & x3))) | (x3 & ((~x1 & ~x4) | (~x2 & ~x8))) | (x1 & ~x3 & ~x8));
endmodule