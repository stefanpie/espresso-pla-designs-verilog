module pla__ti ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    x42, x43, x44, x45, x46,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    x41, x42, x43, x44, x45, x46;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71;
  assign z00 = (x35 & (x44 ? ((x45 & (x46 ? ((~x43 | (~x42 & x43)) & (x19 | (~x19 & x39 & x40))) : (~x43 | (x42 & x43)))) | (~x42 & ~x45 & ~x46)) : (x45 ? ~x46 : (x42 ? ((x43 & (x46 ? ((~x20 | (x20 & x21 & x22)) & ((x18 & x19) | (x39 & x40))) : ((x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))))) | (x11 & x13 & ~x39 & ~x43 & x46 & (x40 | (x19 & ~x40)))) : (x46 & (x43 | (~x43 & (~x21 | ~x22) & (~x18 | ~x19 | (x18 & x19))))))))) | (~x35 & ~x42 & x43 & x44 & x45 & ~x46);
  assign z01 = x35 & (x44 ? ((~x46 & ((x42 & (x43 | (~x43 & x45))) | (~x45 & (~x43 | (~x42 & x43))))) | (~x42 & ~x43 & x45 & x46 & (x19 | (~x19 & x39 & x40)))) : (x45 ? ((x42 & x43 & x46) | (~x43 & ~x46)) : (x42 ? ((x43 & (x46 ? (((~x20 | (x20 & x21 & x22)) & ((x18 & x19) | (x39 & x40))) | (~x20 & ~x36 & (~x18 | ~x19) & (~x39 | ~x40))) : (((x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))) | (~x03 & (~x22 | (~x20 & x21 & x22 & ~x36)) & (~x01 | (x41 & (x05 | x06))))))) | (~x39 & ~x43 & x46 & (((x40 | (x19 & ~x40)) & (~x13 | (x11 & x13))) | (~x19 & ~x40)))) : (x43 | (~x43 & x46 & ((~x22 & (~x18 | ~x19 | (x18 & x19))) | (~x20 & ~x36)))))));
  assign z02 = x35 & (x44 ? ((x45 & x46 & (x19 | (~x19 & x39 & x40)) & (x42 ^ x43)) | (~x46 & (x42 | (~x42 & x43 & ~x45)))) : (x45 ? (x43 ? ((x42 & x46) | (~x19 & ~x42 & ~x46)) : ~x46) : (x42 ? ((x43 & (x46 ? (((~x18 | ~x19) & (~x39 | ~x40)) | (~x20 & ((x18 & x19) | (x39 & x40)))) : (((x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))) | (~x03 & (~x01 | (x41 & (x05 | x06))) & (~x22 | (x21 & x22)))))) | (~x39 & ~x43 & x46 & ((~x19 & ~x40) | (~x13 & (x40 | (x19 & ~x40)))))) : (x43 | (~x43 & x46 & ((~x21 & (~x18 | ~x19)) | ~x20 | (x20 & x21 & x22) | (~x13 & x18 & x19 & ~x22)))))));
  assign z03 = x35 & ((x42 & (x44 ? (x43 ? (~x45 & ~x46) : (x45 & x46 & (x19 | (~x19 & x39 & x40)))) : ((~x45 & ((x46 & ((~x39 & ~x43 & ((~x19 & ~x40) | (~x11 & x13 & (~x19 ^ ~x40)))) | (x20 & x21 & x22 & x43 & ((x18 & x19) | (x39 & x40))))) | (~x11 & ~x22 & x43 & ~x46 & ((~x04 & ~x05 & ~x06) | (x03 & x41))))) | (x43 & x45 & ~x46)))) | (x44 & ((x45 & x46 & (x19 ? (~x42 & x43) : (x40 & (x39 ? (~x42 & x43) : ~x43)))) | (~x42 & ~x43 & ~x46))) | (~x42 & ~x44 & ((x43 & ~x45 & ~x46) | (x19 & ((x43 & x45 & ~x46) | (x18 & ~x21 & ~x43 & ~x45 & x46))))));
  assign z04 = x35 & ((~x44 & (x45 ? (~x46 & (~x43 | (~x18 & x42 & x43))) : ((x46 & ((x19 & ((x18 & ((x20 & x21 & x22 & x42 & x43) | (x13 & ~x22 & ~x42 & ~x43))) | (x42 & ~x43 & ~x39 & ~x40))) | (~x43 & ((~x39 & x40 & x42 & (~x13 | (x13 & (x11 | (~x11 & ~x19))))) | (~x21 & ~x42 & (~x18 | ~x19)))) | (x20 & x21 & x22 & x39 & x40 & x42 & x43))) | (x42 & x43 & ~x46 & ((~x22 & ((~x05 & ~x06 & (x11 | (x04 & ~x11))) | (x11 & (x03 | (x01 & ~x03 & ~x41))) | (~x03 & (~x01 | (x41 & (x05 | x06)))))) | (~x41 & ((x01 & ~x03 & (~x11 | (x21 & x22))) | (x03 & ~x11))) | (x21 & x22 & (x03 | (~x05 & ~x06)))))))) | (x44 & ((x45 & ((x42 & ((~x19 & x39 & x40 & ~x43 & x46) | (x43 & ~x46))) | (x46 & (x19 ? ~x43 : (x40 & ~x42 & (~x43 | (~x39 & x43))))))) | (x42 & ~x43 & ~x46))) | (~x42 & x43 & ~x45 & ~x46));
  assign z05 = x35 & ~x44 & ~x45 & x46 & ((x05 & ((~x06 & (x07 ? (x08 & (x04 ? (~x30 & ~x32) : (~x29 & ~x33))) : (~x08 & (x04 ? (~x30 | ~x32) : (~x29 | ~x33))))) | (x04 & x06 & ((~x30 & (~x08 | (x07 & x08 & ~x33))) | (~x07 & ~x33))))) | (x06 & ((~x05 & ((~x33 & (x04 ? (~x32 & (~x07 | (x07 & x08 & ~x29 & ~x30))) : (~x07 | (x07 & x08 & (~x29 | ~x30))))) | (~x30 & (x04 ? (~x08 & ~x29) : (~x08 | (x07 & x08 & ~x32)))))) | (~x04 & ((~x29 & (~x08 | (x07 & x08 & ~x32))) | (~x07 & ~x32))))));
  assign z06 = x35 & ((~x44 & ((~x45 & (x42 ? (x43 & ((~x46 & (((~x22 | (x21 & x22)) & ((~x05 & ~x06) | (~x03 & (~x01 | (x41 & (x05 | x06)))))) | ((~x07 | x08) & (x04 ? x05 : (x06 | (x05 & ~x06)))) | (x05 & (x07 | ~x08)) | ((x22 ? x21 : x11) & (x03 | ~x41)) | (~x11 & ((x03 & (~x41 | (~x22 & x41))) | (x01 & ~x03 & ~x41) | (~x22 & (~x19 | (~x18 & x19))))) | (~x05 & x06))) | (~x39 & x46 & (x40 | (x18 & ~x19 & ~x40))))) : (~x43 & x46 & (x22 ? x21 : (~x18 | ~x19))))) | (~x40 & x42 & x43 & x45 & x46))) | (x42 & x43 & x44 & ~x45 & ~x46));
  assign z07 = x35 & ((x42 & x43 & x44 & ~x45 & ~x46) | (~x44 & ((~x45 & (x42 ? (x43 ? ((~x46 & (((~x22 | (x21 & x22)) & ((~x05 & ~x06) | (~x03 & (~x01 | (x41 & (x05 | x06)))))) | ((~x07 | x08) & (x04 ? x05 : (x06 | (x05 & ~x06)))) | (x05 & (x07 | ~x08)) | ((x22 ? x21 : x11) & (x03 | ~x41)) | (~x11 & ((x03 & (~x41 | (~x22 & x41))) | (x01 & ~x03 & ~x41) | (~x22 & (~x19 | (~x18 & x19))))) | (~x05 & x06))) | (~x18 & ~x19 & ~x39 & ~x40 & x46)) : x46) : (~x43 & x46 & (x22 ? x21 : (~x18 | ~x19))))) | (x43 & x45 & x46 & ~x39 & x42))));
  assign z08 = x35 & ((x42 & ((~x44 & ((~x45 & ((~x11 & x19 & ((x13 & ~x39 & ~x40 & ~x43 & x46) | (x43 & ~x46 & ~x18 & ~x22))) | (x38 & x43 & x46))) | (x45 & x46 & ~x38 & x43))) | (~x45 & ~x46 & x43 & x44))) | (~x19 & ~x39 & x40 & x44 & x45 & x46));
  assign z09 = x35 & ((~x19 & ~x39 & x40 & x44 & x45 & x46) | (x42 & ((~x45 & ~x46 & x43 & x44) | (~x44 & ((~x45 & ((~x11 & x19 & ((x13 & ~x39 & ~x40 & ~x43 & x46) | (x43 & ~x46 & ~x18 & ~x22))) | (x43 & x46 & x37 & ~x38))) | (~x37 & x43 & x46))))));
  assign z10 = x35 & (x44 ? ((~x46 & (x42 ? (x43 & ~x45) : ((~x43 & x45) | (~x12 & x43 & ~x45)))) | (~x19 & ~x39 & x40 & x45 & x46)) : (x45 ? (~x46 & (~x42 | (x42 & x43))) : (x42 ? ((x43 & (x46 ? (x37 | (~x37 & x38)) : ((x41 & (x05 | x06) & ((x21 & x22) | (x03 & x11 & ~x22))) | (~x04 & ~x05 & ~x06 & (x22 ? x21 : x11)) | (~x11 & ~x22 & (~x19 | (~x18 & x19))) | (x21 & x22 & ~x01 & ~x03)))) | (~x39 & ~x43 & x46 & ((~x19 & ~x40) | (~x11 & x13 & (~x19 ^ ~x40))))) : (~x43 & x46 & (x22 ? x21 : ~x10)))));
  assign z12 = x35 & (x44 ? ((~x19 & ~x39 & x40 & x45 & x46) | (x42 & x43 & ~x45 & ~x46)) : ((~x45 & ((x42 & ((~x11 & ((x13 & ~x39 & ~x43 & x46 & (~x19 ^ ~x40)) | (~x22 & x43 & ~x46 & (~x19 | (~x18 & x19))))) | (x43 & ((~x03 & x21 & x22 & ~x46 & (~x01 | (x41 & (x05 | x06)))) | (x37 & x46))) | (~x40 & ~x43 & x46 & ~x19 & ~x39))) | (x21 & x22 & ~x42 & ~x43 & x46))) | (x45 & ~x46 & ~x42 & x43)));
  assign z13 = x35 & (x44 ? ((~x19 & ~x39 & x40 & x45 & x46) | (x42 & x43 & ~x45 & ~x46)) : ((~x45 & (x42 ? ((~x11 & x19 & ((x13 & ~x39 & ~x40 & ~x43 & x46) | (x43 & ~x46 & ~x18 & ~x22))) | (x43 & ((~x03 & x21 & x22 & ~x46 & (~x01 | (x41 & (x05 | x06)))) | (x38 & x46)))) : (~x43 & x46 & (x22 ? x21 : ~x10)))) | (x45 & ~x46 & x42 & x43)));
  assign z14 = x35 & (x44 ? ((~x19 & ~x39 & x40 & x45 & x46) | (x42 & x43 & ~x45 & ~x46)) : ((x45 & ~x46 & ~x42 & x43) | (~x45 & (x42 ? ((~x11 & ((x13 & ~x39 & ~x43 & x46 & (~x19 ^ ~x40)) | (~x22 & x43 & ~x46 & (~x19 | (~x18 & x19))))) | (~x40 & ~x43 & x46 & ~x19 & ~x39) | (x43 & ((~x03 & x21 & x22 & ~x46 & (~x01 | (x41 & (x05 | x06)))) | (~x37 & x38 & x46)))) : (~x43 & x46 & (x22 ? x21 : ~x10))))));
  assign z15 = x35 & ~x44 & ((x43 & x45 & ~x46) | (~x45 & ((x42 & ((~x19 & ((~x11 & ((x40 & ~x43 & x46 & x13 & ~x39) | (~x22 & x43 & ~x46))) | (~x39 & ~x40 & ~x43 & x46))) | (x43 & x46 & (~x37 ^ ~x38)))) | (~x10 & ~x22 & ~x42 & ~x43 & x46))));
  assign z16 = x35 & (x44 ? ((~x19 & ~x39 & x40 & x45 & x46) | (x42 & x43 & ~x45 & ~x46)) : ((x45 & ~x46 & x42 & x43) | (~x45 & (x42 ? ((~x11 & ((x13 & ~x39 & ~x43 & x46 & (~x19 ^ ~x40)) | (~x22 & x43 & ~x46 & (~x19 | (~x18 & x19))))) | (~x40 & ~x43 & x46 & ~x19 & ~x39) | (x43 & ((~x03 & x21 & x22 & ~x46 & (~x01 | (x41 & (x05 | x06)))) | (x37 & ~x38 & x46)))) : (~x43 & x46 & (x22 ? x21 : ~x10))))));
  assign z17 = x35 & ((~x19 & ~x39 & x40 & x44 & x45 & x46) | (~x45 & ((~x44 & (x42 ? ((x46 & ((~x39 & ~x43 & ((~x19 & ~x40) | (~x11 & x13 & (~x19 ^ ~x40)))) | (x43 & (x37 | (~x37 & x38))))) | (x43 & ~x46 & ((~x11 & ~x22 & (~x19 | (~x18 & x19))) | (~x03 & x21 & x22 & (~x01 | (x41 & (x05 | x06))))))) : (~x43 & x46 & (x22 ? x21 : ~x10)))) | (x42 & x43 & x44 & ~x46))));
  assign z18 = x35 & ~x46 & ((x43 & ((x42 & ~x44 & (x45 | (~x45 & (x22 ? x21 : x11) & ((~x04 & ~x05 & ~x06) | (x03 & x41 & (x05 | x06)))))) | (~x12 & ~x42 & x44 & ~x45))) | (~x42 & x45 & (~x44 | (~x43 & x44))));
  assign z19 = x46 & ~x45 & ~x44 & ~x43 & ~x42 & x35 & ~x10 & ~x22;
  assign z20 = x35 & x46 & ((x26 & x27 & x28 & x44 & x45) | (x23 & x24 & x25 & x42 & ~x43 & ~x44 & ~x45));
  assign z21 = x35 & x46 & ((x28 & x44 & x45 & ~x26 & x27) | (x42 & ~x43 & ~x44 & ~x45 & ~x23 & x24 & x25));
  assign z22 = x35 & x46 & ((x28 & x44 & x45 & x26 & ~x27) | (x42 & ~x43 & ~x44 & ~x45 & x23 & ~x24 & x25));
  assign z23 = x35 & x46 & ((x28 & x44 & x45 & ~x26 & ~x27) | (x42 & ~x43 & ~x44 & ~x45 & ~x23 & ~x24 & x25));
  assign z24 = x35 & x46 & ((x23 & x24 & x25 & x44 & x45) | (x42 & ~x43 & ~x44 & ~x45 & x26 & x27 & x28));
  assign z25 = x35 & x46 & ((x25 & x44 & x45 & ~x23 & x24) | (x42 & ~x43 & ~x44 & ~x45 & ~x26 & x27 & x28));
  assign z26 = x35 & x46 & ((x25 & x44 & x45 & x23 & ~x24) | (x42 & ~x43 & ~x44 & ~x45 & x26 & ~x27 & x28));
  assign z27 = x35 & x46 & ((x25 & x44 & x45 & ~x23 & ~x24) | (x42 & ~x43 & ~x44 & ~x45 & ~x26 & ~x27 & x28));
  assign z28 = x35 & ((x42 & ((~x44 & ((~x09 & ~x46 & (x43 ? (~x45 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))) : x45)) | (~x43 & ~x45 & x46 & ~x27 & ~x28))) | (x44 & x45 & ~x46 & x17 & ~x43))) | (x44 & ((x45 & x46 & ~x24 & ~x25) | (x43 & ~x45 & ~x46 & ~x09 & x12 & ~x42))));
  assign z29 = x35 & (x44 ? (x45 & ((~x27 & ~x28 & x46) | (~x43 & ~x46 & x05 & ~x42))) : ((x42 & ((~x43 & ~x45 & x46 & ~x24 & ~x25) | (x45 & ~x46 & x12 & x43))) | (x43 & x45 & ~x46 & x15 & ~x42)));
  assign z30 = x35 & (x44 ? (x45 & ((x26 & ~x27 & ~x28 & x46) | (~x42 & ~x43 & ~x46 & x04 & x05))) : ((x42 & ((~x43 & ~x45 & x46 & x23 & ~x24 & ~x25) | (x43 & x45 & ~x46 & x11 & x12))) | (x43 & x45 & ~x46 & x14 & x15 & ~x42)));
  assign z31 = x35 & ((x42 & ((~x44 & ((~x09 & ~x46 & (x43 ? (~x45 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))) : x45)) | (~x43 & ~x45 & x46 & x26 & ~x27 & ~x28))) | (x44 & x45 & ~x46 & x16 & x17 & ~x43))) | (x44 & ((x43 & ~x45 & ~x46 & ~x09 & x12 & ~x42) | (x23 & ~x24 & ~x25 & x45 & x46))));
  assign z32 = ~x46 & x45 & x44 & x43 & ~x35 & ~x42;
  assign z33 = x35 & ~x46 & ((x42 & (x43 ? (x44 ? x45 : (~x45 & ((x09 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))) | ((x07 | ~x08) & (x05 ? ~x04 : x06))))) : (x45 & ((x16 & ~x17 & x44) | (x09 & ~x44))))) | (x09 & x12 & ~x42 & x43 & x44 & ~x45));
  assign z34 = x35 & ~x46 & ((x42 & ((x43 & ((~x44 & ~x45 & (((x07 | ~x08) & (x04 ? (x05 | (~x05 & x06 & ~x29)) : (~x05 & x06))) | (x09 & ~x29 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))))) | (~x29 & x44 & x45))) | (~x29 & ~x43 & x45 & ((x16 & ~x17 & x44) | (x09 & ~x44))))) | (x09 & x12 & ~x29 & ~x42 & x43 & x44 & ~x45));
  assign z35 = ~x29 & ~x30 & x35 & ~x46 & ((x09 & ((x42 & ~x44 & (x43 ? (~x45 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))) : x45)) | (x12 & ~x42 & x43 & x44 & ~x45))) | (x16 & ~x17 & x42 & ~x43 & x44 & x45));
  assign z36 = (~x35 & ~x42 & x43 & x44 & x45 & ~x46) | (x35 & (x44 ? (x45 & ((~x26 & x27 & ~x28 & x46) | (~x42 & ~x43 & ~x46 & x04 & ~x05))) : ((x42 & ((~x43 & ~x45 & x46 & ~x23 & x24 & ~x25) | (x43 & x45 & ~x46 & x11 & ~x12))) | (x43 & x45 & ~x46 & x14 & ~x15 & ~x42))));
  assign z37 = x35 & ((x42 & ((~x44 & ((x09 & ~x46 & (x43 ? (~x45 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))) : x45)) | (~x26 & x46 & ((x24 & x43) | (x27 & ~x28 & ~x43 & ~x45))))) | (x44 & x45 & ~x46 & x16 & ~x17 & ~x43))) | (x44 & ((~x23 & x24 & ~x25 & x45 & x46) | (x43 & ~x45 & ~x46 & x09 & x12 & ~x42))));
  assign z38 = x46 & ~x44 & x43 & x42 & x35 & ~x24 & ~x26;
  assign z39 = x35 & ((x44 & ((~x23 & x24 & ~x25 & x45 & x46) | (x43 & ~x45 & ~x46 & x09 & x12 & ~x42))) | (x42 & ((x44 & x45 & ~x46 & x16 & ~x17 & ~x43) | (~x44 & (x43 ? ((x09 & ~x45 & ~x46 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))) | (~x26 & x46 & (~x24 ^ x25))) : ((~x26 & x27 & ~x28 & ~x45 & x46) | (x09 & x45 & ~x46)))))));
  assign z40 = ~x26 & x35 & x42 & x43 & ~x44 & x46 & (x24 ^ x25);
  assign z41 = x35 & ((x44 & ((~x23 & x24 & ~x25 & x45 & x46) | (x43 & ~x45 & ~x46 & x09 & x12 & ~x42))) | (x42 & ((x44 & x45 & ~x46 & x16 & ~x17 & ~x43) | (~x44 & ((x09 & ~x46 & (x43 ? (~x45 & (x22 ? x21 : x11) & (~x41 | (x04 & ~x05 & ~x06))) : x45)) | (~x26 & x46 & (x43 | (x27 & ~x28 & ~x43 & ~x45))))))));
  assign z42 = x35 & x42 & x43 & ~x44 & ~x45 & ~x46 & (~x07 | x08) & ((x06 & (~x04 | ~x05)) | (x04 & x05 & ~x06));
  assign z43 = x35 & x42 & x43 & ~x44 & ~x45 & ~x46 & (~x07 | x08) & ((x06 & (x04 ? (x05 | (~x05 & ~x32)) : ~x05)) | (~x04 & x05 & ~x06));
  assign z45 = x35 & (x44 ? (x45 & ((x26 & x27 & ~x28 & x46) | (~x42 & ~x43 & ~x46 & ~x04 & ~x05))) : ((x42 & ((~x43 & ~x45 & x46 & x23 & x24 & ~x25) | (x43 & x45 & ~x46 & ~x11 & ~x12))) | (x43 & x45 & ~x46 & ~x14 & ~x15 & ~x42)));
  assign z46 = x35 & ((x46 & ((x24 & ((x26 & x42 & x43 & ~x44) | (x44 & x45 & x23 & ~x25))) | (x42 & ~x43 & ~x44 & ~x45 & x26 & x27 & ~x28))) | (~x16 & ~x17 & x42 & x45 & ~x46 & ~x43 & x44));
  assign z47 = x46 & ~x44 & x43 & x42 & x35 & ~x24 & x26;
  assign z48 = x35 & ((~x16 & ~x17 & x42 & x45 & ~x46 & ~x43 & x44) | (x46 & ((x24 & ((x44 & x45 & x23 & ~x25) | (x25 & x26 & x42 & x43 & ~x44))) | (x26 & x42 & ~x44 & ((x27 & ~x28 & ~x43 & ~x45) | (~x24 & ~x25 & x43))))));
  assign z49 = x26 & x35 & x42 & x43 & ~x44 & x46 & (x24 ^ x25);
  assign z50 = x35 & ((x42 & ((x26 & ~x44 & x46 & (x43 | (x27 & ~x28 & ~x43 & ~x45))) | (x44 & x45 & ~x46 & ~x16 & ~x17 & ~x43))) | (x44 & x45 & x46 & x23 & x24 & ~x25));
  assign z51 = (~x35 & ~x42 & x43 & x44 & x45 & ~x46) | (x35 & (x44 ? (~x46 & (x42 ? (~x43 & x45) : (x43 & ~x45))) : ((x42 & x43 & (x46 | (~x45 & ~x46 & (x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))))) | (~x43 & ((x45 & ~x46) | (~x10 & ~x22 & ~x42 & ~x45 & x46))))));
  assign z52 = (~x35 & ~x42 & x43 & x44 & x45 & ~x46) | (x35 & (x44 ? (~x46 & (x42 ? (~x43 & x45) : (x43 & ~x45))) : ((~x45 & (x42 ? (x43 & (x46 ? (((~x20 | (x20 & x21 & x22)) & ((x18 & x19) | (x39 & x40))) | ((~x18 | ~x19) & (~x39 | ~x40)) | x28 | ~x37 | x38 | (~x39 & x40) | (x37 & ~x38)) : ((x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))))) : (~x43 & x46 & ((x18 & x19 & (~x21 | (x13 & ~x22))) | ~x20 | (x20 & x21 & x22) | (~x10 & ~x22))))) | (~x43 & x45 & ~x46))));
  assign z54 = ~x46 & ((x35 & ((x42 & (x43 ? (~x44 & ~x45 & (x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))) : (x44 & x45))) | (~x42 & x43 & x44 & ~x45) | (~x43 & ~x44 & x45))) | (~x35 & ~x42 & x43 & x44 & x45));
  assign z55 = ~x46 & ~x45 & x44 & ~x43 & x35 & x42;
  assign z56 = ~x46 & ~x45 & x44 & ~x43 & x35 & ~x42;
  assign z57 = ~x46 & ~x45 & x44 & ~x43 & x35 & x42;
  assign z58 = x46 & ~x44 & x43 & x42 & ~x28 & x35;
  assign z59 = x46 & ~x44 & x43 & x42 & x28 & x35;
  assign z60 = x46 & ~x44 & x43 & x42 & x35 & ~x27 & ~x28;
  assign z62 = x35 & ~x43 & ~x45 & ((~x10 & ~x22 & ~x42 & ~x44 & x46) | (x42 & x44 & ~x46));
  assign z63 = x35 & ((x27 & ~x28 & x42 & x43 & ~x44 & x46) | (~x42 & ~x43 & x44 & ~x45 & ~x46));
  assign z64 = x35 & x42 & ~x45 & ((~x44 & x46 & x28 & x43) | (~x43 & x44 & ~x46));
  assign z65 = x46 & ~x45 & ~x44 & x43 & x42 & x35 & ~x20 & x28;
  assign z66 = x35 & x42 & ~x45 & ((~x43 & x44 & ~x46) | (x43 & ~x44 & x46 & x20 & x28));
  assign z68 = x46 & ~x45 & ~x44 & x43 & x42 & x35 & x27 & x28;
  assign z69 = x46 & ~x45 & ~x44 & x43 & x42 & x35 & ~x27 & x28;
  assign z70 = (~x35 & ~x42 & x43 & x44 & x45 & ~x46) | (x35 & ((~x46 & ((x42 & (x43 ? (~x44 & ~x45 & (x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))) : (x44 & x45))) | (~x42 & x43 & x44 & ~x45) | (~x43 & ~x44 & x45))) | (~x10 & ~x22 & ~x42 & ~x45 & x46 & ~x43 & ~x44)));
  assign z71 = ~x46 & ((x35 & ((x42 & (x43 ? (~x44 & ~x45 & (x22 ? x21 : x11) & (x03 | (~x05 & ~x06) | (x01 & ~x03 & ~x41))) : (x44 & x45))) | (~x42 & x43 & x44 & ~x45) | (~x43 & ~x44 & x45))) | (~x35 & ~x42 & x43 & x44 & x45));
  assign z11 = 1'b0;
  assign z44 = 1'b0;
  assign z53 = 1'b0;
  assign z61 = 1'b0;
  assign z67 = 1'b0;
endmodule