module pla__prom1 ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39;
  assign z00 = (x2 & ((x4 & ((x1 & ((~x0 & ((x5 & ((x3 & ~x6 & (~x7 | (x7 & ~x8))) | (x6 & (~x7 | (x7 & x8))))) | (~x3 & ((~x5 & (~x7 | (x7 & x8))) | (x6 & x7 & ~x8))))) | (~x3 & ((x5 & (~x6 | (x0 & x6 & x7))) | (x0 & (x7 ? ~x5 : x6)))) | (x0 & x3 & ~x5 & x6 & ~x7))) | (~x1 & ((x5 & (x0 ? (x6 & ((x3 & (~x7 ^ x8)) | (~x7 & x8))) : ((~x6 & ~x7) | (~x3 & x7 & ~x8)))) | (x0 & ((~x3 & (~x6 | (x6 & x7 & x8))) | (~x5 & x6 & (~x7 | (x3 & x7))))))) | (x3 & (x0 ? (~x5 & ~x6) : (x5 & x7 & (x6 ^ x8)))))) | (x5 & ((~x4 & ((~x0 & (x6 ? x3 : ~x1)) | (x3 & ((x0 & x6 & (x7 | (x1 & ~x7))) | (x1 & ~x6))) | (x0 & ~x1 & ((x6 & ~x7) | (~x3 & (x8 ? x7 : ~x6)))))) | (~x1 & (x0 ? ((x3 & ~x6) | (x7 & ~x8 & ~x3 & x6)) : (~x3 & x6 & (~x7 | (x7 & x8))))))) | (~x4 & ((~x5 & (x0 ? (~x1 | (x1 & x3)) : x3)) | (x1 & ~x3))) | (~x0 & ~x1 & ~x3 & ~x5))) | (x3 & ((x4 & (x5 ? ((~x6 & ((x1 & ~x2) | (x7 & ~x8 & ~x0 & ~x1))) | (~x1 & (((~x7 | (x7 & x8)) & (x0 ? ~x2 : x6)) | (x7 & ~x8 & x0 & x6))) | (x1 & ~x2 & x6 & (x0 ? (~x8 | (x7 & x8)) : x7))) : (~x0 | (x0 & ~x2)))) | (~x2 & (x0 ? ~x4 : ((~x4 & ((~x5 & (x1 ? ~x7 : (~x6 & x8))) | (~x8 & (x1 ? (x6 ? x7 : x5) : (~x6 & x7))) | (~x1 & x6 & (~x7 | (x7 & x8))) | (x1 & x7 & x8))) | (x5 & ((x6 & (x1 ? ~x7 : (x7 & ~x8))) | (~x1 & ~x6 & (~x7 | (x7 & x8)))))))))) | (~x2 & ~x3);
  assign z01 = x0 ? (x2 & ~x3 & ~x5 & ((x1 & ~x4 & ~x7 & (x6 ^ x8)) | (~x1 & x4 & ~x6 & x7 & ~x8))) : ((~x1 & ((~x5 & ~x6 & ((x2 & ((~x3 & x8 & (~x4 | (x4 & ~x7))) | (~x4 & x7 & ~x8))) | (~x2 & x3 & ~x4 & x7 & x8))) | (~x2 & x3 & x4 & x5 & x6 & (~x7 ^ ~x8)))) | (x1 & x2 & ~x3 & x4 & ~x7 & x8 & ~x5 & x6));
  assign z02 = (x0 & ((~x1 & ((~x2 & ((~x4 & (~x3 | (x7 & x8 & x3 & x5))) | (x4 & ((x3 & x5 & (x6 ? x8 : x7)) | (~x5 & ((x6 & x7 & x8) | (~x3 & (~x7 | (x7 & ~x8))))))) | (x3 & (x5 ? (~x6 & ~x7) : (~x6 | (x6 & ~x7)))))) | (x2 & ((x3 & ((~x7 & ((~x4 & (x8 ? x6 : ~x5)) | (~x6 & x8 & x4 & x5))) | (x4 & ((~x5 & x6 & x8) | (x7 & ~x8 & x5 & ~x6))))) | (~x5 & ((~x3 & ~x4) | (~x7 & ~x8 & x4 & x6))) | (x5 & ((~x3 & ((~x4 & x7 & x8) | (x6 & ~x7 & ~x8))) | (~x7 & (x4 ? (x6 ^ ~x8) : ~x6)))) | (~x3 & x4 & (x6 ? (x7 & x8) : (~x7 ^ ~x8))))) | (x6 & ~x8 & ((x7 & ((x4 & x5) | (x3 & (~x4 | (x4 & ~x5))))) | (x3 & x5 & ~x7))))) | (x5 & ((x1 & (x2 ? (x3 ? (~x4 & ((x7 & ~x8) | (x6 & (~x7 ^ x8)))) : (x4 & (~x6 ^ x7))) : ((x3 & ~x7 & ((x6 & x8) | (x4 & (~x6 | (x6 & ~x8))))) | (~x4 & ((~x6 & ~x8) | (~x3 & x6 & x8)))))) | (~x3 & x4 & ((~x2 & (~x6 | (x6 & ~x7))) | (x7 & x8 & x2 & ~x6))))) | (x1 & ((~x2 & ((~x5 & (x3 ? (x7 ? (x4 | (~x4 & ~x8)) : ~x6) : (x4 | (~x4 & ~x7)))) | (~x4 & ((x7 & x8 & ~x3 & ~x6) | (~x7 & ~x8 & x3 & x6))))) | (~x5 & ((x6 & ((x2 & x7 & (~x3 | (x3 & ~x4))) | (x3 & x4 & ~x7))) | (x2 & ~x3 & x4 & ~x6))) | (x2 & ~x3 & (x4 ? (x6 & ~x7) : ~x6)))) | (x2 & x3 & x4 & ~x5 & ~x6))) | (~x0 & ((x6 & ((x1 & (x3 ? ((x4 & ((x2 & ~x8 & (~x5 | (x5 & ~x7))) | (~x2 & x5 & ~x7) | (~x5 & x7 & x8))) | (~x2 & ~x4 & (~x7 | (x5 & x7 & x8)))) : ((x4 & ~x5) | (~x2 & ~x4 & x8)))) | (~x1 & ((x5 & (x7 ? ((~x2 & (~x3 | (x3 & x8))) | (~x8 & (x3 ? x4 : x2))) : (x2 ? (x4 ^ x8) : x4))) | (x2 & ~x5 & ((x4 & ~x7) | (~x3 & ~x4 & x8))) | (~x2 & ~x4 & ~x7))) | (x2 & x5 & ((x3 & ~x7 & (x4 ^ ~x8)) | (x4 & x7 & x8))) | (x7 & ~x8 & x3 & ~x4))) | (~x6 & ((x1 & ((x2 & x4 & (~x5 | (~x7 & x8 & x3 & x5))) | (~x3 & ((~x2 & ~x5) | (~x4 & x5 & x7))) | (~x2 & x3 & ((x5 & ~x7) | (~x4 & (x8 ? x7 : ~x5)))))) | (x5 & ((~x1 & (x2 ? ((x7 & (x8 ? ~x3 : x4)) | (x3 & ~x7 & x8)) : (~x3 | (x3 & x4)))) | (x2 & x3 & (x4 ? (~x7 ^ x8) : (x7 & ~x8))))) | (~x1 & (x2 ? (~x5 & ~x7) : (x3 & ~x4))))) | (~x5 & (x2 ? (x1 ? (~x3 & ~x4) : (x7 & (x4 | (~x3 & ~x4 & ~x8)))) : ((x4 & (~x1 | (x1 & x3 & (~x7 | (x7 & ~x8))))) | (~x1 & ~x3 & ~x4 & x7)))) | (~x3 & x5 & ((x1 & ((x4 & ~x7) | (x2 & (x4 ? (x7 & ~x8) : ~x7)))) | (~x1 & x2 & ~x4 & ~x7 & ~x8))))) | (x3 & ((x2 & ~x4 & ((x8 & ((x5 & (x1 ? (~x6 ^ ~x7) : (x6 & x7))) | (~x1 & ~x5 & x7))) | (x1 & (x5 ? (~x6 & ~x7) : (~x6 | (x6 & ~x7)))))) | (x1 & ~x2 & x4 & x5 & x7 & (~x6 | (x6 & ~x8))))) | (x1 & x5 & x6 & x7 & (x2 ? (~x3 & ~x4) : (x8 ? x4 : ~x3)));
  assign z03 = (x2 & ((~x4 & (x3 ? ((x7 & ((x0 & (x1 ? (x5 ? ~x8 : x6) : (x8 ? (~x5 | (x5 & ~x6)) : x6))) | (~x0 & ((x1 & ((x6 & ~x8) | (x5 & ~x6 & x8))) | (x5 & ~x6 & ~x8))) | (x6 & x8 & ~x1 & x5))) | (~x0 & ((~x1 & x8 & (x5 ? ~x7 : x6)) | (~x5 & ~x6) | (~x7 & ~x8 & x5 & x6))) | (x0 & (x1 ? (x5 ? (~x7 & (~x6 | (x6 & ~x8))) : ~x6) : ((x6 & ~x7) | (~x5 & ~x6 & ~x8)))) | (x1 & x6 & ~x7 & (~x5 | (x5 & x8)))) : ((~x6 & ((x0 & x1) | (~x0 & ~x1 & x5 & ~x8))) | (x7 & (x0 ? (x1 ? (x6 & ~x8) : (x5 & x8)) : (x1 ? (x5 & x8) : (~x5 & ~x8)))) | (x1 & (x0 ? (x6 & x8) : ~x5)) | (~x1 & (x0 ? (~x5 | (x5 & ~x7)) : (~x5 & ~x7))) | (x6 & ~x7 & ~x0 & x5)))) | (x4 & ((x0 & ((x1 & ((~x3 & (~x5 | (x5 & (~x6 ^ x7)))) | (x6 & ~x7 & x3 & ~x5))) | (~x1 & ((x5 & ((~x8 & (x3 ? (~x6 ^ ~x7) : ~x6)) | (x6 & ~x7 & x8))) | (x6 & x7 & x8) | (~x3 & ~x7 & (x6 ^ x8)))) | (~x3 & x5 & ~x6 & x7 & x8))) | (x5 & ((x1 & ((~x0 & ~x8 & (x3 ? (x6 & ~x7) : (~x6 & x7))) | (~x3 & x6 & ~x7))) | (~x0 & ((~x1 & (x6 ? (~x7 & ~x8) : (~x7 | (x7 & ~x8)))) | (x6 & x7 & x8) | (x3 & (x6 ? (~x7 ^ ~x8) : (x7 & x8))))))) | (~x0 & ~x5 & (~x6 | (x6 & ((~x1 & (~x7 | (x7 & ~x8))) | (x3 & (x8 ? x7 : x1)))))))) | (~x0 & ~x3 & ((x7 & ((~x1 & x8 & (~x5 ^ ~x6)) | (x5 & x6 & ~x8))) | (~x6 & ~x7 & x1 & x5))))) | (~x2 & ((x5 & ((~x3 & ((~x1 & ((x0 & x4 & ~x6) | (x7 & ~x8 & ~x0 & ~x4))) | (~x6 & ((~x4 & (x0 ? (x1 & ~x8) : x8)) | (x0 & x1 & x7 & (x8 | (x4 & ~x8))))) | (x6 & ((x0 & ((x4 & ~x7) | (x1 & x7 & ~x8))) | (x7 & x8 & ~x0 & x1))) | (x4 & ~x7 & ~x0 & x1))) | ((~x6 | (x6 & ~x7)) & ((~x0 & ~x1 & x4) | (x3 & ~x4 & x0 & x1))) | (x4 & ((x7 & ((~x0 & ((x6 & ~x8) | (x1 & ~x6 & x8))) | (x0 & (x1 ? ((x6 & x8) | (x3 & (x6 ^ x8))) : (x3 & ~x6))) | (~x6 & ~x8 & x1 & x3))) | (x0 & ((x1 & ~x6 & ~x7) | (x6 & x8 & ~x1 & x3))) | (x6 & ~x7 & x1 & x3))) | (~x1 & ((x0 & x3 & ((~x4 & x7 & x8) | (x6 & ~x7 & ~x8))) | (x7 & x8 & ~x0 & x6))))) | (~x4 & (x0 ? (x1 ? (x3 ? (~x5 & (~x7 | (x7 & ~x8))) : (x6 & (~x7 | (x7 & x8)))) : (~x3 | (x3 & ~x5))) : ((~x5 & (x1 ? (x3 ? (~x6 & ~x8) : (x6 & x8)) : (~x3 & x7))) | (~x1 & (x6 ? ~x7 : x3)) | (x1 & ((x6 & x7 & ~x8) | (x3 & (x7 ? x8 : x6))))))) | (~x5 & ((x4 & (x0 ? (x1 ? x6 : ((x6 & x7 & x8) | (~x3 & ~x7))) : (~x1 | (x1 & x3 & (~x7 | (x7 & ~x8)))))) | (x1 & ~x3 & ~x6))) | (~x0 & x1 & x3 & x7 & x8 & x4 & x6))) | (~x0 & ((x3 & ((~x6 & ~x7 & x1 & x5) | (x6 & x7 & ~x8 & ~x1 & ~x4))) | (x1 & ~x3 & ((x4 & ~x5 & x6) | (~x6 & x7 & ~x8 & ~x4 & x5))))) | (x0 & ((x3 & ((x5 & ((~x1 & ~x6 & ~x7) | (x6 & x7 & x8 & x1 & ~x4))) | (x4 & ~x5 & (~x6 | (~x1 & x6 & (~x7 | (x7 & ~x8))))))) | (~x1 & x4 & x7 & ~x8 & (x5 ? x6 : ~x3))));
  assign z04 = (x4 & ((~x0 & ((~x2 & ((~x3 & ((~x5 & (x7 ? x8 : ~x1)) | (~x1 & (x6 ? (x7 & ~x8) : x5)) | (x1 & ~x6 & ~x8))) | (x8 & ((x3 & ~x5 & (x6 ? x7 : x1)) | (x1 & x5 & (x7 | (x6 & ~x7))))) | (x1 & ((~x5 & x6 & ~x7) | (~x6 & ~x8 & x3 & x5))) | (~x1 & ((~x7 & ~x8 & x5 & x6) | (x3 & ~x5 & (~x6 | (x6 & ~x8))))))) | (x2 & ((x5 & ((x8 & ((x6 & (~x7 | (x3 & x7))) | (x1 & (x3 ? (~x6 & ~x7) : x7)))) | (~x6 & (x1 ? (~x3 & ~x7) : (x7 & ~x8))))) | (x1 & x3 & ((x7 & ~x8) | (~x5 & ~x7 & x8))) | (~x3 & ((~x1 & ~x7 & (x8 ? ~x5 : x6)) | (x7 & x8 & ~x5 & x6))) | (x7 & ~x8 & ~x1 & ~x5))) | (~x1 & x3 & x5 & (x6 ? (x7 & ~x8) : ~x7)) | (x6 & x7 & ~x8 & x1 & ~x3 & ~x5))) | (x0 & ((x2 & ((~x7 & ((x1 & x3 & ~x5) | (~x3 & x5 & x6))) | (~x1 & ((~x8 & ((x3 & (x5 ? ~x6 : x7)) | (x5 & x6 & x7))) | (~x3 & (~x5 | (x5 & ~x6))))) | (x1 & ((~x3 & ((~x5 & (~x6 | (x6 & x7))) | (x7 & x8 & x5 & x6))) | (~x6 & x7 & ~x8 & x3 & ~x5))))) | (x6 & ((~x2 & (((x3 | (~x3 & x8)) & (x1 ? ~x5 : ~x7)) | (x7 & ~x8 & ~x1 & ~x5) | (x1 & ((~x3 & x7 & ~x8) | (x5 & ((~x7 & ~x8) | (x3 & (~x7 ^ ~x8)))))))) | (~x5 & x7 & x8 & ~x1 & x3))) | (~x6 & ((x1 & ((~x2 & ~x5) | (~x3 & x5 & ~x8))) | (x5 & ((~x1 & x7 & (x8 ? x3 : ~x2)) | (~x2 & x3 & ~x7))) | (~x3 & ~x7 & ~x1 & ~x2))) | (~x2 & ~x3 & x7 & x8 & (~x1 ^ x5)))) | (~x1 & ((x2 & x3 & ~x7 & (~x5 | (x5 & x6 & ~x8))) | (x6 & x7 & x8 & ~x2 & x5))) | (~x5 & x6 & ~x7 & x1 & x2 & ~x3))) | (~x4 & ((~x0 & ((x3 & ((~x1 & ((x5 & (x2 ? ~x7 : (~x6 & x8))) | (x6 & x7 & ~x8) | (~x2 & ((x6 & ~x7) | (~x5 & ~x6 & ~x8))))) | (x5 & (x6 ^ ~x8) & (x2 ? x1 : x7)) | (x2 & ((~x5 & ~x6) | (~x7 & ~x8 & x1 & x6))) | (x1 & ~x5 & x7 & (x8 ? x6 : ~x2)))) | (x1 & ((x5 & ((~x3 & ~x6) | (~x2 & x6 & ~x7))) | (~x3 & ((~x2 & x7 & (x8 ? ~x5 : x6)) | (x6 & ~x8 & x2 & ~x5))) | (~x2 & ~x5 & ~x7))) | (~x3 & ((~x1 & (~x2 | (x2 & ~x6 & (x8 ? ~x5 : x7)))) | (x7 & x8 & x2 & x6))))) | (x5 & ((~x3 & ((x0 & ~x1 & ~x6) | (x6 & ~x7 & x1 & x2))) | (x0 & ((~x6 & ((x1 & x2) | (~x1 & ~x2 & x3 & ~x8))) | (x3 & ((x6 & ((x1 & (~x7 | (x2 & x7 & x8))) | (x2 & x7 & ~x8))) | (~x1 & (x2 ? (~x7 & ~x8) : (x7 & x8))))) | (~x1 & ~x2 & x6 & (~x7 | (x7 & ~x8))))) | (x3 & ~x6 & ((x1 & ~x2 & ~x7) | (x7 & x8 & ~x1 & x2))))) | (x0 & ((~x5 & ((x7 & ((x1 & (x2 ? (~x3 & ~x8) : (x3 & x8))) | (~x3 & x8 & ~x1 & x2))) | (~x7 & (x1 ? (x2 ^ x3) : (~x2 & ~x3))) | (x2 & x3) | (~x1 & ~x8 & (x2 ? (~x3 & ~x6) : (x3 & x6))))) | (~x3 & (x1 ? (~x2 | (x7 & x8 & x2 & x6)) : (x6 & x7 & (x2 ^ x8)))) | (x6 & x7 & ~x8 & x1 & ~x2 & x3))) | (~x1 & ((x6 & ~x7 & x2 & ~x3) | (~x2 & x3 & ~x5 & x7 & x8))))) | (~x6 & (x0 ? (~x2 & x3 & (x1 ? (x5 & x7) : (~x5 & ~x7))) : (x2 & ~x3 & (x1 ? ~x5 : (x5 & (~x7 | (x7 & x8))))))) | (x5 & x6 & ((x7 & ((~x8 & ((~x0 & ((x2 & ~x3) | (x1 & ~x2 & x3))) | (x2 & ~x3 & x0 & x1))) | (x0 & x8 & (x1 ? (~x2 & x3) : (x2 & ~x3))))) | (x0 & ~x1 & x2 & x3 & x8)));
  assign z05 = (x3 & ((x5 & ((~x4 & ((~x0 & (x2 ? (~x6 & ((x7 & x8) | (x1 & ~x8) | (~x1 & ~x7))) : ((x6 & (~x7 | (x7 & x8))) | (~x1 & (x8 ? ~x6 : x7))))) | (x0 & ((x1 & (x2 ? (x7 ? ~x8 : ~x6) : (~x6 | (x6 & ~x7)))) | (x2 & ((x6 & ~x7) | (~x1 & x7 & x8))) | (~x1 & ~x8 & (~x6 | (x6 & x7))))) | (x6 & x7 & x8 & x1 & x2))) | ((x0 ? (x4 & x7) : ~x7) & ((x1 & ~x2 & ~x6) | (x6 & ~x8 & ~x1 & x2))) | (x4 & ((x6 & ((x8 & ((~x7 & (x0 ? (~x1 ^ ~x2) : ~x1)) | (~x0 & (x2 ? x7 : x1)))) | (x7 & ~x8 & (x0 ? (x1 & ~x2) : ~x1)))) | (x2 & ~x8 & (x0 ? (~x1 & ~x7) : (x1 & x7))) | (~x6 & (x0 ? ((~x2 & ~x7) | (~x1 & x7 & x8)) : ((~x1 & ~x7) | (~x2 & x7 & x8)))))) | (x6 & ((~x2 & ((x0 & (x1 ? (x7 & x8) : ~x7)) | (x7 & ~x8 & ~x0 & x1))) | (~x0 & x1 & x2 & ~x7))))) | (~x1 & ((~x5 & ((x4 & ((x6 & (x0 ? ~x7 : (~x2 & ~x8))) | (~x0 & (x2 ? ~x7 : ~x6)) | (x0 & (x2 ? (x7 ? ~x8 : ~x6) : (x7 & x8))))) | (~x2 & (x0 ? ((~x6 & ~x7) | (~x4 & x6 & ~x8)) : (~x4 & (x6 | (~x6 & ~x8))))))) | (x7 & ((x0 & x8 & (x2 ? (x4 & x6) : ~x4)) | (~x4 & x6 & ~x8 & ~x0 & x2))) | (x6 & ~x7 & x8 & ~x0 & x2 & ~x4))) | (~x5 & ((x1 & (x4 ? ((~x6 & ((~x0 & (x8 ? ~x2 : x7)) | (x2 & (~x7 | (x0 & x7))))) | (x0 & x6 & (~x2 | (x2 & ~x7)))) : ((x7 & x8 & ~x0 & x6) | (x0 & ~x2 & (~x7 | (x7 & x8)))))) | (~x0 & ((x2 & ~x4 & ~x6) | (x6 & x7 & x8 & ~x2 & x4))) | (x0 & x2 & ~x4))) | (x1 & ~x2 & ~x4 & x7 & ~x8 & (~x0 ^ x6)))) | (x2 & ((~x0 & ((~x7 & ((~x1 & ~x3 & x6) | (x5 & ~x6 & x1 & x4))) | (~x5 & ((~x1 & ((x4 & x7 & ~x8) | (~x3 & ~x6 & x8))) | (~x3 & ((x1 & ~x6) | (x7 & x8 & x4 & x6))) | (x1 & x6 & ~x8 & (~x4 | (x4 & x7))))) | (x7 & ((~x3 & ((~x1 & ~x6 & (x8 ? x5 : ~x4)) | (x6 & (x8 ? ~x4 : x5)))) | (~x1 & x4 & x5 & ~x6 & ~x8))))) | (~x3 & ((x0 & ((x7 & ((~x6 & ((~x1 & ~x4) | (x5 & x8 & x1 & x4))) | (~x1 & (x4 ? x5 : (x6 & ~x8))) | (x1 & ((~x4 & (~x8 | (x6 & x8))) | (x6 & ~x8 & x4 & x5))))) | (x4 & (~x5 | (x5 & x6 & ~x7))) | (~x4 & ~x7 & (x1 | (~x1 & x6))))) | (x5 & ((~x1 & ~x6 & ~x7) | (x6 & x7 & x8 & x1 & x4))))))) | (~x2 & ((x4 & ((x0 & ((~x6 & ((x1 & ~x5) | (x7 & ~x8 & ~x1 & x5))) | (~x1 & ((~x3 & x5 & ~x7) | (x7 & ~x8 & ~x5 & x6))) | (x1 & ((x5 & ((x6 & ~x7 & ~x8) | (~x3 & x7 & x8))) | (~x3 & x6 & (x8 ? ~x5 : x7)))))) | (~x1 & ((~x3 & ((~x5 & ~x7) | (~x0 & (x5 ? ~x6 : (x6 & x7))))) | (x5 & x6 & ((x7 & x8) | (~x0 & ~x7 & ~x8))))) | (~x0 & x1 & ~x3 & ~x6 & ~x8))) | (~x3 & ((x5 & ((x0 & ~x4) | (x6 & x7 & x8 & ~x0 & x1))) | (~x5 & ((x1 & (x0 ? ~x4 : (x7 & x8))) | (x0 & ~x1 & (x7 ? x8 : ~x4)))) | (~x0 & ((~x1 & ~x4) | (x7 & ~x8 & x1 & x6))))) | (~x0 & x1 & ~x4 & ~x5 & ~x7))) | (x1 & ((~x0 & ((x4 & ((~x5 & x6 & ~x7) | (~x3 & x5 & ~x6 & x7 & x8))) | (~x3 & x5 & (x6 ? ~x7 : ~x4)))) | (x5 & ~x6 & ~x8 & x0 & ~x3 & x4)));
  assign z06 = (x5 & ((~x0 & ((x1 & ((x6 & ((~x2 & x8 & (x3 ? ~x4 : x7)) | (x3 & (x4 ? ~x7 : (x7 & ~x8))) | (x4 & ~x7 & x2 & ~x3))) | (x4 & ((~x6 & (x2 ? (x3 ? ~x7 : ~x8) : x3)) | (~x2 & ~x3 & ~x7))) | (~x4 & ((~x2 & ~x6) | (~x7 & x8 & x2 & ~x3))))) | (~x1 & ((~x2 & ((~x4 & (x3 ? (x8 ? x7 : ~x6) : (x7 & ~x8))) | (~x3 & ~x7 & (~x6 | (x6 & ~x8))) | (~x6 & x8 & x3 & x4))) | (x6 & ((~x3 & x7 & x8) | (x4 & ~x7 & (x8 | (x3 & ~x8))))) | (~x6 & ~x7 & x2 & x4))) | (x2 & ((x3 & ((~x4 & (~x6 | (x6 & x7 & x8))) | (x7 & ~x8 & x4 & ~x6))) | (x4 & x7 & (x6 ^ x8)))) | (x4 & x7 & ((~x2 & ~x3 & ~x6) | (x3 & x6 & x8))))) | (x2 & ((x0 & (x1 ? (x3 ? (~x4 & (x7 ? (~x8 | (x6 & x8)) : ~x6)) : (~x6 | (x6 & (x4 ? (x8 | (x7 & ~x8)) : ~x7)))) : ((x6 & x7 & x8) | (x4 & (x7 ? (x6 ^ x8) : ((~x3 & ~x8) | (x6 & (x8 | (x3 & ~x8))))))))) | (~x1 & ((~x3 & ~x6 & (x8 ? ~x4 : x7)) | (~x4 & x6 & ~x7))) | (x1 & x3 & ~x4 & x6 & ~x7))) | (x0 & ((x3 & ((~x4 & ((~x1 & ~x6) | (x6 & ~x7 & x1 & ~x2))) | (~x2 & ((x1 & ((x6 & x7 & x8) | (x4 & ~x6 & ~x7))) | (x7 & ~x8 & x4 & ~x6) | (~x1 & x6 & ~x7))) | (~x6 & ~x7 & ~x1 & x4))) | (x1 & ~x2 & x4 & x6 & ~x7))) | (~x2 & x6 & x7 & ~x8 & (x1 ? x4 : x3)))) | (x1 & ((~x3 & (((x2 ? ~x5 : ~x4) & (x0 | (~x0 & x6 & ~x7))) | (~x2 & ((~x6 & ((x0 & x4) | (~x5 & ~x8 & ~x0 & ~x4))) | (x6 & ((x7 & ~x8 & ~x0 & ~x4) | (x0 & x4 & (x8 ? x7 : ~x5)))) | (~x5 & x7 & x8 & ~x0 & ~x4))) | (~x0 & x2 & ((~x5 & ((~x6 & x8) | (x4 & x7 & ~x8))) | (x7 & (x8 ? x6 : ~x4)))))) | (x3 & ((~x5 & (x4 ? ((x0 & (~x6 | (~x2 & x6 & x7))) | (x2 & x6 & (~x7 | (~x0 & x7 & ~x8)))) : (x2 ? (x0 ? (x8 ? x7 : ~x6) : (~x6 | (x6 & x7))) : (~x0 | (x0 & x6 & x8))))) | (x0 & ~x2 & ~x4 & (~x6 | (x6 & x7 & ~x8))))) | (x4 & ~x5 & ~x0 & ~x2))) | (~x1 & ((~x5 & ((x4 & (x3 ? (x0 ? (x2 ? (x6 & (x8 | (x7 & ~x8))) : (x8 ? ~x6 : x7)) : ((x6 & (~x7 | (x7 & ~x8))) | (~x2 & ~x6 & ~x8))) : (x2 | (~x0 & ~x2 & (~x7 | (x7 & x8)))))) | (~x4 & ((x0 & ((~x2 & x3) | (x7 & x8 & x2 & ~x3))) | (~x0 & (~x2 | (x2 & ((x7 & x8) | (x3 & ~x6 & ~x8))))) | (x2 & ~x3 & ~x7))) | (x3 & ~x6 & x0 & x2))) | (~x2 & ((x0 & (~x3 | (x6 & x7 & x8 & x3 & x4))) | (x6 & x7 & ~x8 & ~x0 & ~x3 & x4))) | (x6 & x7 & ~x8 & x2 & ~x4))) | (x3 & ~x5 & ((x2 & ((~x4 & x6 & ~x7) | (~x0 & x4 & (~x6 | (x6 & x7 & x8))))) | (x0 & ~x2 & x4 & x6 & ~x7)));
  assign z07 = (x2 & ((x6 & ((x4 & ((x0 & (x1 ? (~x3 & ((~x5 & ~x7) | (x7 & ~x8) | (x5 & x8))) : ((x3 & (x5 ? (~x7 & ~x8) : (x8 | (x7 & ~x8)))) | (x5 & (~x7 ^ ~x8))))) | (~x5 & (x3 ? ((x1 & ~x7) | (~x0 & x7 & (x8 | (x1 & ~x8)))) : ((x1 & x7 & x8) | (~x0 & ~x7)))) | (~x0 & x5 & (x7 ? ~x8 : (x8 | (x3 & ~x8)))))) | (~x4 & ((~x1 & (x0 ? ((~x3 & x7 & ~x8) | (x5 & ~x7)) : (~x7 & (x8 ? ~x3 : x5)))) | (x7 & ((~x0 & ~x8 & (~x3 | (x3 & ~x5))) | (x3 & x8 & (x5 | (x1 & ~x5))))) | (~x7 & ((x3 & ~x5) | (x1 & x5 & (x3 | (x0 & ~x3))))))) | (x5 & x7 & x8 & x0 & ~x1 & ~x3))) | (x0 & ((~x6 & (x5 ? ((x3 & (x1 ? (~x4 & ~x7) : (x4 & x8))) | (~x3 & (x1 ? (~x4 | (x4 & (~x7 | (x7 & ~x8)))) : (x8 ? ~x4 : x7))) | (~x7 & ~x8 & ~x1 & x4)) : (x1 ? (x3 ? ((x4 & (~x7 | (x7 & ~x8))) | (x7 & x8) | (~x4 & ~x8)) : x4) : (x3 & x4)))) | (~x4 & (x1 ? ((~x3 & ~x5) | (x7 & ~x8 & x3 & x5)) : (~x3 & ~x5 & (~x7 | (x7 & x8))))) | (x4 & ~x5 & ~x1 & ~x3))) | (~x0 & ((~x3 & (x5 ? ((x1 & ~x8 & (x7 ? ~x6 : x4)) | (~x4 & ~x6 & x8)) : ((~x1 & ~x6 & ~x7) | (x4 & (x1 ? (x8 ? ~x6 : x7) : x7))))) | (x3 & ~x6 & ((x1 & ((~x4 & ~x5) | (x7 & ~x8 & x4 & x5))) | (~x4 & (x5 | (~x1 & ~x5 & ~x8))) | (x4 & (~x5 | (x5 & (~x7 | (x7 & x8))))))) | (~x5 & x7 & x8 & ~x1 & ~x4))) | (x1 & ~x3 & x4 & x7 & x8 & x5 & ~x6))) | (~x0 & ((~x3 & ((~x6 & ((~x1 & x4 & x5) | (x1 & ~x2 & ~x4 & ~x5 & ~x8))) | (~x4 & ((~x2 & ((x7 & ~x8 & x1 & x6) | (~x1 & x5 & (~x7 | (x7 & ~x8))))) | (x1 & ((x6 & ~x7) | (~x5 & x7 & x8))))) | (x6 & ((x5 & x7 & x8) | (~x2 & x4 & ((~x1 & x7 & ~x8) | (x5 & ~x7))))) | (~x1 & ~x2 & x4 & ~x5 & (~x7 | (x7 & x8))))) | (x3 & ((~x2 & ((~x4 & (x1 ? (~x5 | (x5 & x6 & x8)) : (x5 & (x8 ? x7 : ~x6)))) | (~x1 & ((x4 & ~x6 & (x5 ^ ~x8)) | (x7 & ~x8 & x5 & x6))))) | (x4 & ((x7 & ((x5 & x6 & x8) | (~x1 & ~x8 & (~x5 ^ ~x6)))) | (x6 & ~x7 & ~x1 & ~x5))) | (x6 & x7 & ~x8 & x1 & ~x4 & x5))) | (~x2 & (x1 ? (x5 ? ~x6 : x4) : (~x4 & ~x5))))) | (x0 & ((~x2 & ((x1 & ((x6 & ((~x5 & (x3 ? (~x4 & x8) : (x4 & ~x8))) | (~x3 & x4 & (x7 ? x8 : x5)) | (x3 & ((x5 & x7 & x8) | (~x4 & (x7 ? ~x8 : x5)))))) | (~x3 & (~x4 | (x4 & ~x6))) | (x3 & ~x6 & (~x4 | (x4 & x5 & (~x7 | (x7 & ~x8))))))) | (~x1 & (~x3 | (x3 & (x4 ? (x5 & (~x7 | (x7 & ~x8))) : (x6 & ~x7))))) | (x3 & x4 & ~x5))) | (~x1 & x3 & ((~x4 & (~x6 | (x6 & x7 & ~x8))) | (x6 & x7 & x8 & x4 & x5))))) | (x1 & ~x2 & x4 & x5 & x6 & (x7 ? ~x8 : x3));
  assign z08 = (x0 & ((~x1 & ((x2 & (x3 ? ((~x5 & (~x6 | (x4 & x6 & x8))) | (x6 & x7 & ~x8) | (x5 & ((x4 & (x6 ? (~x7 & ~x8) : (x7 & x8))) | (~x7 & (~x6 | (x6 & x8)))))) : ((x6 & (x4 ? (~x7 | (x5 & x7)) : (x5 & x8))) | (x5 & ~x6) | (~x4 & ~x5 & ~x7)))) | (~x3 & ((~x2 & (x4 ? (x5 ? (x8 ? ~x6 : x7) : ~x6) : ((x6 & ~x7) | (~x5 & ~x6 & ~x8)))) | (~x4 & x7 & (x8 ? ~x5 : x6)))) | (~x2 & ((x4 & ((~x5 & ((x6 & ~x7) | (x3 & x7 & ~x8))) | (x3 & ~x6 & (~x7 | (x5 & x7))))) | (x5 & ((~x4 & ~x6) | (x3 & x6 & ~x7))))) | (x6 & x7 & x8 & x3 & x4 & x5))) | (x6 & (x2 ? ((x1 & ((x3 & ((~x4 & x7) | (~x7 & ~x8 & x4 & ~x5))) | (x5 & ((~x4 & ~x7) | (~x3 & x4 & (x8 | (x7 & ~x8))))))) | (x3 & ~x4 & ~x5 & ~x7)) : ((x4 & ((x7 & ((~x5 & x8) | (x1 & ((x5 & ~x8) | (x3 & (x5 ^ ~x8)))))) | (x1 & ~x7 & ((~x3 & ~x8) | (x5 & (x8 | (x3 & ~x8))))))) | (~x3 & x5 & ((x7 & x8) | (x1 & ~x4 & ~x8)))))) | (x1 & ((x4 & ((~x6 & (x2 ? (x3 ? (~x5 & x7) : x5) : (x3 ? (~x5 | (x5 & x7 & ~x8)) : (~x5 & x8)))) | (~x3 & ~x5 & (x2 | (~x2 & x7 & ~x8))))) | (~x4 & (x3 ? (x2 ? (~x6 & (~x5 | (x5 & x7))) : x5) : ~x5)) | (x5 & ~x6 & ~x2 & ~x3))))) | (~x0 & ((x5 & ((x1 & ((~x3 & ((x6 & x7 & ~x8) | (~x6 & x8 & ~x2 & x4))) | (x3 & ((x6 & ((x4 & ((~x7 & x8) | (x2 & (~x7 ^ x8)))) | (~x2 & (x8 ? x7 : ~x4)))) | (x7 & x8 & (x4 ? ~x6 : x2)))) | (~x2 & (x4 ? (~x8 & (~x6 ^ ~x7)) : ~x6)))) | (~x1 & ((x2 & (((~x6 ^ ~x7) & (x8 ? x4 : ~x3)) | (x6 & x7 & x8) | (~x3 & ~x6 & ~x7))) | (~x2 & (x3 ? ((x8 & (x7 | (x6 & ~x7))) | (x4 & ~x6 & ~x8)) : (~x6 | (x6 & x7)))) | (x3 & ~x7 & (x4 ? (x6 & ~x8) : ~x6)))) | (x2 & x3 & x4 & (x7 ? ~x8 : ~x6)))) | (~x5 & ((x4 & ((x1 & ((~x2 & (~x3 | (x3 & ~x6 & ~x8))) | (x7 & ~x8 & x2 & x6))) | (x3 & (((~x6 | (x6 & x8)) & (x7 ? x2 : ~x1)) | (~x2 & x7 & x8) | (x6 & ~x8 & (x7 ? ~x1 : x2)))))) | (~x4 & ((x2 & ((x3 & ((x7 & x8) | (x1 & ~x6 & ~x8))) | (~x1 & ~x6 & ~x8))) | (x1 & ~x3 & (x8 ? ~x6 : x7)))) | (~x1 & ~x3 & (~x2 | (x2 & x6 & ~x7))))) | (x2 & ((~x4 & ((x3 & x6 & ~x7) | (x7 & ((~x1 & ((x6 & ~x8) | (~x3 & ~x6 & x8))) | (x6 & ~x8 & x1 & x3))))) | (x1 & ~x3 & x4 & ((x6 & ~x7) | (x7 & x8) | (~x6 & ~x8))))) | (x1 & x6 & ((~x3 & ~x4 & (~x7 | (x7 & x8))) | (~x2 & x3 & x4 & x7 & ~x8))))) | (x2 & (x4 ? (~x5 & (x1 ? (x3 & ~x7 & (~x6 | (x6 & x8))) : (~x3 & (~x6 | (x6 & x7))))) : (x5 & ~x6 & (x1 ? (~x3 | (x3 & ~x7)) : (x3 & x7))))) | (~x2 & ((x3 & ((x1 & x4 & ~x7 & (~x5 ^ ~x6)) | (~x4 & ~x5) | (x6 & x7 & ~x8 & ~x1 & x5))) | (x5 & x6 & ~x7 & ~x1 & ~x3 & x4)));
  assign z09 = (x6 & ((x0 & ((~x2 & ((~x3 & ((~x4 & (x1 ? (x5 & ~x8) : ~x7)) | (x1 & ((x5 & x7 & x8) | (x4 & ~x7 & ~x8))))) | (~x7 & ((x4 & (x1 ? (x5 & (x8 | (x3 & ~x8))) : ~x5)) | (~x1 & x3 & x5))) | (x4 & x7 & ((x5 & ~x8) | (x1 & ((~x5 & x8) | (x3 & (x5 ^ ~x8)))))))) | (x1 & ((x3 & ((x2 & ~x4 & (x5 ? (~x8 | (x7 & x8)) : x7)) | (x4 & ~x5 & ~x7))) | (x2 & ~x3 & x5 & (x4 ? (x8 | (x7 & ~x8)) : ~x7)))) | (~x1 & (x3 ? ((~x4 & ((x2 & ~x5 & ~x7) | (x5 & x7 & ~x8))) | (x2 & ((x4 & (~x5 ^ ~x8)) | (~x5 & x7 & ~x8) | (x5 & ~x7 & x8))) | (x7 & x8 & x4 & x5)) : ((x4 & ((~x5 & x7 & x8) | (x2 & (~x7 | (x7 & ~x8))))) | (x7 & (x8 ? x5 : ~x4))))))) | (~x0 & ((x5 & (x1 ? ((x3 & ((x4 & ((x7 & ~x8) | (~x7 & x8) | (x2 & (~x7 ^ x8)))) | (~x4 & ~x7 & ~x8) | (~x2 & x7 & x8))) | (~x3 & (x7 ? ~x8 : ~x4)) | (~x7 & ~x8 & ~x2 & x4)) : ((~x7 & ((x2 & (x8 ? x4 : ~x3)) | (x3 & (x8 ? ~x2 : x4)))) | (x2 & x7 & x8) | (~x2 & ((~x3 & ~x4 & x8) | (x7 & (~x8 | (x4 & x8)))))))) | (x2 & ((~x5 & ((x4 & ((x1 & (x8 ? x3 : x7)) | (~x1 & (x8 ? x7 : ~x3)) | (x3 & ~x7 & ~x8))) | (~x3 & (x1 ? (~x4 & ~x8) : (~x7 & x8))))) | (x1 & ((x7 & ~x8 & x3 & ~x4) | (~x3 & x4 & ~x7))) | (~x1 & ~x4 & (x7 ? ~x8 : x3)))) | (x7 & ((x1 & ~x3 & ((~x4 & x8) | (~x2 & x4 & ~x5))) | (~x1 & x3 & x4 & ~x5 & ~x8))) | (~x5 & ~x7 & x8 & ~x1 & x3 & x4))) | (~x7 & ((x1 & x2 & x3 & ~x4 & (~x5 | (x5 & x8))) | (~x1 & ~x2 & ~x3 & x4 & x5))))) | (~x6 & ((x1 & ((~x0 & ((~x2 & (x4 ? ((x5 & (~x7 ^ ~x8)) | (x3 & x7 & x8)) : ((x5 & x7 & x8) | (~x3 & (x8 ? ~x7 : x5))))) | (x2 & (x3 ? (x4 ? (x5 & (x8 | (x7 & ~x8))) : (~x5 & ~x8)) : (x4 & ~x8))) | (x3 & x4 & x5 & ~x7 & ~x8))) | (x3 & ((x0 & ((x4 & (x2 ? (~x5 & x7) : (~x5 | (x5 & ~x7)))) | (x2 & ~x4 & (~x5 | (x5 & x7))))) | (~x5 & ~x7 & x2 & x4))) | (~x3 & ((x5 & ((x2 & ~x4) | (x0 & (~x2 | (x2 & x4 & x7))))) | (x0 & ~x2 & x4 & ~x5 & x8))))) | (~x1 & ((~x0 & ((x5 & ((~x2 & (~x3 | (x3 & x4 & ~x8))) | (x2 & ~x3 & ~x7) | (x7 & x8 & x3 & x4))) | (x2 & ~x4 & ((~x5 & ~x8) | (~x3 & x7 & x8))) | (x3 & x4 & ~x5 & ~x7))) | (x0 & (x2 ? (x3 ? (~x5 | (x7 & x8 & x4 & x5)) : (~x4 & x5)) : (x4 ? (~x5 | (x5 & x8)) : (x5 | (~x3 & ~x5 & ~x8))))) | (x2 & ((x5 & (x3 ? (~x4 ^ ~x7) : (x4 & x7))) | (~x3 & x4 & ~x5))))) | (x3 & ((x5 & (x0 ? ((x2 & ~x4 & ~x7) | (x7 & ~x8 & ~x2 & x4)) : (~x4 & ~x7))) | (~x0 & x2 & x4 & ~x5 & x7))) | (x0 & x2 & ~x3 & x4 & x5 & ~x7))) | (~x5 & (x3 ? ((~x2 & ~x4) | (~x0 & ((~x2 & x4 & (x1 ? ~x8 : (x7 & x8))) | (x7 & x8 & x2 & ~x4)))) : (x0 ? ((~x4 & (x1 | (~x1 & (x7 ? x8 : x2)))) | (x1 & x4 & (x2 | (~x2 & x7 & ~x8)))) : (~x2 & (~x1 | (x1 & (x4 ? ~x7 : (x7 & ~x8)))))))) | (~x0 & x7 & ((x3 & x5 & ((~x4 & (x1 ? (x2 ^ ~x8) : (~x2 & x8))) | (x4 & ~x8 & ~x1 & x2))) | (x1 & x2 & ~x3 & x4 & x8))) | (x0 & x1 & ~x2 & x3 & ~x4 & x5);
  assign z10 = (x4 & ((~x0 & ((~x2 & (x8 ? ((~x7 & ((x1 & ((x5 & x6) | (x3 & ~x5 & ~x6))) | (x5 & ~x6 & ~x1 & x3))) | (~x1 & x3 & x5 & x6 & x7)) : ((x1 & ((x3 & (x5 ? (x6 & ~x7) : (~x6 & x7))) | (~x6 & x7 & ~x3 & x5))) | (~x5 & x6 & ~x7 & ~x1 & ~x3)))) | (x2 & ((~x8 & ((x1 & ((~x3 & ~x5 & x7) | (~x6 & ~x7 & x3 & x5))) | (~x6 & ~x7 & ~x1 & ~x3))) | (~x1 & x8 & ((x3 & ~x5 & x7) | (x5 & ((~x6 & x7) | (~x3 & x6 & ~x7))))))) | (~x6 & x7 & ~x8 & ~x1 & ~x3 & ~x5))) | (x0 & (x6 ? (x1 ? ((x2 & ((~x3 & x5 & x7) | (~x7 & ~x8 & x3 & ~x5))) | (x5 & x8 & ((~x3 & ~x7) | (~x2 & x3 & x7)))) : ((~x3 & ((x2 & ((~x7 & ~x8) | (~x5 & x7 & x8))) | (x7 & ((~x5 & ~x8) | (~x2 & x5 & x8))))) | (x7 & ~x8 & x3 & x5) | (~x2 & ~x7 & ((x5 & ~x8) | (x3 & ~x5 & x8))))) : ((x7 & ((~x2 & x3 & ((x5 & x8) | (~x1 & ~x5 & ~x8))) | (~x1 & ~x3 & x8 & (~x5 | (x2 & x5))))) | (x2 & ~x3 & ~x5 & ~x7 & (~x1 | (x1 & ~x8)))))) | (x1 & x2 & ~x3 & ~x6 & x8 & (~x5 ^ x7)))) | (~x4 & ((x2 & (x6 ? (x0 ? ((x5 & ((~x1 & x7 & (x3 ^ x8)) | (~x7 & ~x8 & x1 & x3))) | (x1 & ~x5 & (x7 ? x8 : x3))) : ((~x3 & ((x1 & (x5 ? (x7 & ~x8) : (~x7 & x8))) | (~x7 & ~x8 & ~x1 & ~x5))) | (~x1 & x7 & (x5 ? x8 : x3)))) : ((x5 & ((x7 & (x0 ? ((~x3 & ~x8) | (~x1 & x3 & x8)) : (x1 ? x3 : ~x8))) | (x0 & ~x7 & (~x1 ^ x3)))) | (x0 & ~x5 & (x1 ? (x3 & ~x8) : (x7 & x8)))))) | (~x2 & ((x3 & (x8 ? ((x1 & ~x5 & (x0 ? x7 : ~x6)) | (x0 & ~x1 & x7 & (~x6 | (x5 & x6)))) : ((~x5 & (x0 ? (~x1 & (~x6 | (x6 & x7))) : (x7 | (x1 & x6 & ~x7)))) | (~x1 & x5 & ~x6 & (~x7 | (x0 & x7)))))) | (x0 & ((x1 & ~x3 & (x5 ? (x7 & (x6 ^ ~x8)) : (~x7 & x8))) | (x6 & x7 & x8 & ~x1 & ~x5))))) | (~x0 & x3 & ((~x6 & ~x7 & ~x1 & ~x5) | (x6 & x7 & x8 & x1 & x5))))) | (~x1 & ((~x3 & ((~x7 & ((x0 & ~x2 & (x5 ? x8 : (~x6 & ~x8))) | (x5 & ~x6 & x8 & ~x0 & x2))) | (~x6 & x7 & x8 & ~x0 & x2 & ~x5))) | (x7 & x8 & ~x5 & x6 & ~x0 & ~x2 & x3))) | (~x2 & ~x3 & x0 & x1 & ~x7 & x8 & x5 & ~x6);
  assign z11 = (x2 & (x7 ? (x1 ? ((~x5 & (x0 ? (~x4 & ((~x6 & x8) | (x3 & x6 & ~x8))) : (~x3 & ~x8 & (x6 | (x4 & ~x6))))) | (x0 & ~x4 & x5 & ~x6 & (~x8 | (x3 & x8)))) : ((x0 & ((~x8 & ((~x3 & (x4 ? (~x5 & x6) : x5)) | (x3 & x4 & x5 & x6))) | (x6 & x8 & ~x4 & x5))) | (~x0 & ((x8 & ((x3 & (x4 ? ~x5 : x6)) | (x4 & x5 & ~x6))) | (x3 & ~x4 & x5 & ~x6 & ~x8))) | (~x6 & x8 & ~x3 & ~x5))) : ((x0 & ((~x3 & ((x5 & ((~x1 & (x4 ? (x6 & ~x8) : ~x6)) | (~x6 & x8 & x1 & ~x4))) | (~x6 & ~x8 & x4 & ~x5))) | (x1 & x3 & ((~x6 & ~x8 & x4 & ~x5) | (~x4 & (x5 ? (x6 & ~x8) : (~x6 & x8))))))) | (~x3 & ((~x5 & ((~x0 & ~x4 & (x1 ? x6 : (~x6 & ~x8))) | (~x6 & x8 & x1 & x4))) | (~x0 & ~x1 & x5 & ~x6 & (x8 | (x4 & ~x8)))))))) | (~x2 & ((~x6 & ((~x0 & ((~x8 & ((~x1 & (x3 ? (x5 & x7) : (x4 & ~x5))) | (x4 & x5 & ((x3 & ~x7) | (x1 & ~x3 & x7))))) | (x3 & ~x4 & ~x5 & ~x7) | (x1 & ((x3 & ~x5 & x7 & (~x4 | (x4 & x8))) | (~x7 & x8 & ~x3 & x4))))) | (~x5 & ~x7 & x8 & ~x1 & x3 & x4) | (x0 & ((x7 & ((~x1 & x3 & ~x8 & (~x4 | (x4 & ~x5))) | (x1 & ~x3 & x4 & ~x5 & x8))) | (x1 & ~x3 & ~x7 & (x4 ? (~x5 & ~x8) : x8)))))) | (~x0 & ((x6 & ((~x8 & ((x1 & (x3 ? (~x5 & x7) : (x4 & ~x7))) | (x4 & ~x5 & ~x1 & x3))) | (x5 & x7 & x8 & ~x1 & x3))) | (x1 & ~x3 & ~x4 & ~x5 & x7 & ~x8))) | (x0 & x4 & ((x5 & ((x1 & x8 & (~x3 ^ x7)) | (x6 & ~x8 & ~x1 & x3))) | (~x1 & x6 & (x3 ? (~x7 & x8) : x7)))))) | (~x0 & x4 & x5 & x6 & ~x7 & (x1 ? (x3 & ~x8) : (~x3 & x8)));
  assign z12 = (~x7 & (x4 ? ((~x1 & ((~x3 & ((x0 & x5 & (x2 ? (x6 & x8) : (~x6 & ~x8))) | (~x5 & ~x6 & ~x0 & x2))) | (~x2 & x3 & ((~x0 & x8 & (~x5 | (x5 & x6))) | (x6 & ~x8 & x0 & ~x5))))) | (~x0 & x1 & ((~x8 & ((x2 & x6 & (~x3 ^ ~x5)) | (~x5 & ~x6 & ~x2 & ~x3))) | (~x2 & x3 & x5 & ~x6 & x8)))) : (x1 ? ((~x5 & (x0 ? ((~x2 & x3 & x6 & x8) | (~x6 & ~x8 & x2 & ~x3)) : ((~x6 & x8 & x2 & x3) | (x6 & ~x8 & ~x2 & ~x3)))) | (~x0 & ~x3 & x5 & (x2 ? (x6 & x8) : (~x6 & ~x8)))) : ((x3 & ((x5 & (x0 ? (x2 ? (x6 & ~x8) : (~x6 & x8)) : (~x2 & x8))) | (~x0 & x2 & ~x5 & x6 & ~x8))) | (x2 & ((~x5 & x6 & x8 & x0 & ~x3) | (~x6 & ~x8 & ~x0 & x5))))))) | (x7 & ((~x1 & (x6 ? ((x5 & ((~x0 & ((~x2 & ~x4 & x8) | (x2 & ~x3 & x4 & ~x8))) | (x0 & ~x2 & ~x3 & ~x4 & x8))) | (~x0 & ~x2 & x3 & ~x4 & ~x8)) : ((x8 & ((~x0 & (x2 ? (x3 & ~x4) : (x4 & ~x5))) | (x5 & ((x0 & x2 & ~x3) | (~x2 & x3 & x4))))) | (~x3 & ~x8 & (x0 ? (x5 & (x2 ^ ~x4)) : (x2 & ~x5)))))) | (~x0 & x1 & ((x6 & ((x2 & ~x5 & (x3 ? (~x4 & ~x8) : (x4 & x8))) | (~x2 & ~x3 & ~x4 & x5 & x8))) | (x2 & ~x3 & ~x5 & ~x6 & x8))))) | (~x1 & ~x3 & x8 & ((~x0 & x2 & x6 & (~x4 ^ ~x5)) | (x0 & ~x2 & ~x4 & ~x5 & ~x6)));
  assign z13 = (~x6 & ((~x3 & ((~x5 & (x7 ? ((~x0 & x2 & (x1 ? x8 : (~x4 & ~x8))) | (~x2 & ~x4 & x8 & x0 & ~x1)) : ((x1 & ~x8 & (x0 ? (x2 & ~x4) : (~x2 & x4))) | (x0 & ~x1 & (x2 ? (x4 & x8) : ~x4))))) | (x0 & ((x5 & ((x4 & (x1 ? (x2 ? (x7 & x8) : (~x7 & ~x8)) : (x2 ? (x7 & ~x8) : (~x7 & x8)))) | (~x1 & ~x4 & x7 & (x2 ^ ~x8)))) | (~x1 & ~x2 & x4 & ~x7 & ~x8))) | (x5 & ~x7 & ~x8 & x1 & ~x2 & ~x4))) | (x3 & (x0 ? (~x4 & ((x2 & ((x1 & (x5 ? ~x7 : (x7 & ~x8))) | (x7 & x8 & ~x1 & ~x5))) | (~x1 & ~x2 & (x8 ? x5 : ~x7)))) : ((x8 & ((x7 & ((~x1 & (x2 ? ~x4 : (x4 & x5))) | (x1 & x2 & ~x4 & x5))) | (x1 & ~x7 & (x2 ? (~x4 & ~x5) : (x4 & x5))))) | (x1 & x4 & ~x8 & (x2 ? (x5 & ~x7) : (~x5 & x7)))))) | (~x0 & ~x1 & ((~x5 & x7 & x8 & ~x2 & x4) | (x2 & ~x4 & x5 & ~x7 & ~x8))))) | (x6 & (x0 ? (x2 ? ((~x4 & ((~x5 & ((x1 & (x3 ? (~x7 & ~x8) : (x7 & x8))) | (~x7 & x8 & ~x1 & ~x3))) | (x5 & ~x8 & ~x1 & x3))) | (~x3 & x4 & ((~x1 & ~x5 & (~x7 ^ x8)) | (x5 & ((~x7 & x8) | (x1 & x7 & ~x8)))))) : ((~x4 & x8 & (x1 ? ((~x5 & ~x7) | (~x3 & x5 & x7)) : (x5 & (~x3 | (x3 & x7))))) | (~x1 & x4 & ~x7 & ~x8 & (~x3 ^ ~x5)))) : (x2 ? ((~x8 & (x1 ? ((x3 & ~x5 & (~x4 ^ ~x7)) | (~x3 & x4 & x5 & ~x7)) : ((x3 & ~x4 & ~x5) | (~x3 & x4 & x5 & x7)))) | (~x3 & x8 & (x4 ? (~x5 & x7) : (x5 & ~x7)))) : ((~x1 & ((x3 & ((~x7 & x8 & x4 & ~x5) | (x7 & ~x8 & ~x4 & x5))) | (~x7 & x8 & x4 & x5))) | (~x3 & ~x4 & ((x5 & x7 & x8) | (~x7 & ~x8 & x1 & ~x5))))))) | (~x0 & ~x1 & x8 & ((~x2 & x3 & ~x4 & (x5 ^ x7)) | (x2 & ~x3 & x4 & ~x5 & ~x7)));
  assign z14 = (x5 & (x1 ? ((~x0 & (x4 ? (x2 ? ((x7 & x8 & ~x3 & ~x6) | (~x7 & ~x8 & x3 & x6)) : (~x7 & ((x6 & x8) | (x3 & ~x6 & ~x8)))) : (x6 & x7 & ((x3 & x8) | (x2 & ~x3 & ~x8))))) | (x2 & ((~x4 & ~x6 & ((x3 & x7 & ~x8) | (x0 & x8 & (~x3 ^ x7)))) | (x6 & x7 & x8 & x0 & ~x3 & x4))) | (x0 & ~x2 & ~x3 & ~x4 & ~x6 & ~x8)) : (x0 ? ((~x4 & ((x2 & x7 & (x3 ? x8 : (x6 & ~x8))) | (~x2 & ~x3 & ~x6 & ~x7 & x8))) | (~x2 & x4 & x6 & ((~x3 & x7 & ~x8) | (~x7 & x8)))) : (~x6 & ((~x2 & x3 & (x4 ? (~x7 | (x7 & ~x8)) : ~x8)) | (~x4 & x7 & ~x8 & x2 & ~x3)))))) | (~x5 & (x2 ? ((~x4 & (x0 ? (x1 & ((~x6 & x7 & x8) | (x3 & (x6 ? (x8 | (x7 & ~x8)) : ~x7)))) : ((~x1 & ~x7 & (x3 ? ~x6 : ~x8)) | (x6 & ~x8 & x1 & ~x3)))) | (x4 & ~x7 & ~x8 & x0 & x1 & x3)) : (x0 ? ((x7 & ((~x1 & x6 & (x3 ? (~x4 & ~x8) : x8)) | (x8 & (x3 ? ~x4 : (x4 & ~x6))))) | (~x1 & x3 & x4 & ~x6 & ~x7 & x8)) : ((~x8 & ((x4 & ((~x1 & (x3 ? x6 : ~x7)) | (x6 & x7 & x1 & x3))) | (x1 & ~x4 & (x3 ^ x7)))) | (x3 & ((~x6 & x8 & x1 & x4) | (~x1 & x7 & (x4 ? (x6 & x8) : ~x6)))))))) | (x1 & ~x2 & ~x3 & x4 & ~x7 & (x0 ? (~x6 & ~x8) : (x6 ^ x8)));
  assign z15 = (~x2 & ((~x1 & ((x3 & (x0 ? ((~x6 & x8 & x4 & x5) | (~x4 & ~x8 & (x5 ? (~x6 & ~x7) : (x6 & x7)))) : (x4 & (x5 ? (~x6 & ~x7) : (x6 ? (~x8 | (x7 & x8)) : x8))))) | (x7 & ((~x0 & ~x6 & ((x4 & ~x5 & ~x8) | (~x3 & ~x4 & x5 & x8))) | (~x5 & x6 & x8 & x0 & ~x3 & ~x4))) | (~x3 & x5 & ((x0 & x4 & ~x7 & (~x6 | (x6 & x8))) | (x6 & ~x8 & ~x0 & ~x4))))) | (x1 & (x0 ? (x4 ? (x3 ? (x5 & x7 & (x8 | (x6 & ~x8))) : (~x5 & (x6 ? (~x7 & x8) : ~x8))) : (x6 & ((x3 & ~x5 & (~x7 ^ x8)) | (~x7 & x8 & ~x3 & x5)))) : ((~x3 & ((x4 & x5 & (x6 ? x8 : (~x7 & ~x8))) | (~x6 & ~x7 & ~x4 & ~x5))) | (x3 & x4 & ~x5 & ~x6 & ~x7 & x8)))) | (x0 & ~x3 & ~x5 & ((~x7 & x8 & ~x4 & ~x6) | (x7 & ~x8 & x4 & x6))) | (x5 & x6 & ~x7 & ~x0 & x3 & ~x4))) | (x2 & ((~x3 & ((~x8 & (x1 ? ((x6 & ((x0 & x5 & (~x4 ^ ~x7)) | (~x5 & x7 & ~x0 & x4))) | (~x6 & ~x7 & ~x0 & ~x5)) : ((~x4 & x5 & ~x7 & (x6 | (x0 & ~x6))) | (x6 & x7 & ~x0 & x4)))) | (x8 & ((x5 & ((x0 & ((~x6 & ~x7 & ~x1 & x4) | (~x4 & x6 & x7))) | (x6 & x7 & x1 & x4))) | (~x0 & ((~x1 & ~x5 & x6 & (~x4 ^ ~x7)) | (~x6 & ~x7 & x1 & x4))))) | (~x5 & ~x6 & x7 & x0 & ~x1 & ~x4))) | (~x4 & ((x3 & ((~x6 & ((~x0 & ~x8 & (x1 ? x7 : (~x5 & ~x7))) | (x1 & x8 & ((~x5 & ~x7) | (x0 & x5 & x7))))) | (x0 & ((~x5 & ((x1 & ((x7 & ~x8) | (x6 & ~x7 & x8))) | (x7 & x8 & ~x1 & x6))) | (~x7 & ~x8 & x1 & x5))))) | (~x6 & ~x7 & x8 & ~x0 & ~x1 & ~x5))) | (x0 & ~x1 & x3 & x5 & ((x6 & ~x7 & ~x8) | (x4 & ~x6 & x7))))) | (x0 & ~x1 & x3 & ((~x7 & x8 & x4 & ~x5) | (x6 & ((x4 & ~x8 & (~x5 ^ x7)) | (x7 & x8 & ~x4 & x5)))));
  assign z16 = (~x4 & ((x2 & ((x7 & ((~x8 & ((~x6 & (x0 ? (x5 ? x1 : x3) : (~x1 & ~x3))) | (~x0 & x6 & ((~x3 & x5) | (~x1 & x3 & ~x5))))) | (~x5 & ((x1 & (x0 ? (x8 & (~x3 | (x3 & ~x6))) : (~x3 & x6))) | (~x6 & x8 & ~x1 & x3))))) | (~x7 & (x0 ? ((x3 & (x1 ? (x5 ? (~x6 | (x6 & ~x8)) : (~x8 | (x6 & x8))) : (~x5 & ~x6))) | (~x6 & x8 & ~x3 & x5)) : (~x3 & (x5 ? (x6 ? x1 : ~x8) : (x6 & ~x8))))) | (~x0 & x1 & ~x3 & ~x6 & x8))) | (~x2 & ((~x1 & ((x3 & (x7 ? (x0 ? ((~x6 & x8) | (~x5 & x6 & ~x8)) : (x5 ? ~x8 : x6)) : ((~x6 & ~x8) | (~x0 & x5 & x8)))) | (x0 & ~x3 & x5 & ((~x6 & x7 & ~x8) | (~x7 & (x8 | (x6 & ~x8))))))) | (x1 & ((x6 & (x0 ? (~x3 & (x5 ? (x7 & ~x8) : (~x7 & x8))) : (x3 & ~x5 & (~x7 ^ ~x8)))) | (~x0 & x3 & ~x6 & (x5 ? (~x7 & x8) : ~x8)))) | (x6 & x7 & x8 & x0 & ~x3 & x5))) | (x7 & x8 & ~x5 & x6 & x0 & x1 & x3))) | (~x1 & ((x7 & ((x3 & ((~x2 & ((~x0 & x8 & ((x4 & ~x5 & ~x6) | (x5 & x6))) | (x5 & ~x8 & x0 & x4))) | (x0 & x2 & x5 & (x6 ^ x8)))) | (x4 & ((~x3 & ((x0 & ((~x5 & x6 & x8) | (x2 & x5 & ~x8))) | (~x6 & x8 & x2 & x5))) | (~x0 & ~x2 & ~x5 & x6 & ~x8))))) | (~x3 & ((x4 & ((x2 & ((x0 & x6 & (x5 ? ~x7 : ~x8)) | (~x7 & x8 & ~x5 & ~x6))) | (~x0 & ~x2 & ~x5 & (x6 ? ~x7 : x8)))) | (~x6 & ~x7 & ~x8 & x0 & ~x2 & ~x5))) | (x0 & x6 & ~x7 & ((~x2 & x3 & x4 & x5) | (x2 & ~x5 & x8))))) | (x4 & ((x0 & ((x5 & ((x6 & x7 & x8 & x2 & ~x3) | (x1 & ~x2 & x3 & ~x6 & ~x7 & ~x8))) | (x1 & ((x7 & ((~x2 & ~x8 & (x6 ? ~x5 : x3)) | (~x3 & ~x5 & x8 & (~x6 | (x2 & x6))))) | (~x5 & ~x7 & ((x3 & x6 & ~x8) | (x2 & (x3 ? (~x6 & ~x8) : x8)))))))) | (~x0 & ~x3 & ~x5 & (((x6 ^ ~x8) & ((x1 & ~x2 & ~x7) | (x2 & x7))) | (x1 & x6 & ~x8 & (x7 | (x2 & ~x7))))) | (x1 & ~x2 & x3 & ~x7 & x8 & x5 & x6))) | (x2 & ~x3 & x0 & x1 & ~x7 & ~x8 & ~x5 & ~x6);
  assign z17 = (x1 & ((~x2 & ((x5 & (x0 ? ((~x4 & x7 & ((~x6 & ~x8) | (x3 & (x8 | (x6 & ~x8))))) | (~x3 & x8 & (~x6 | (x4 & x6)))) : ((x4 & (x3 ? (~x6 & ~x7) : (x7 & ~x8))) | (x3 & ((x6 & ~x7 & ~x8) | (~x4 & ~x6 & x7))) | (~x3 & ~x4 & (x6 ? (x7 & x8) : (~x7 & ~x8)))))) | (~x5 & ((~x4 & (x0 ? ((x3 & (~x6 ^ ~x7)) | (x7 & x8 & ~x3 & x6)) : (x3 ? (~x6 & x8) : (x7 & ~x8)))) | (~x0 & x3 & x4 & ~x8 & (~x6 | (x6 & x7))))) | (~x3 & ~x7 & ((~x0 & (x6 ^ x8)) | (x6 & ~x8 & x0 & ~x4))))) | (x2 & ((x4 & ((x5 & ((~x3 & ((~x6 & x7) | (x0 & x6 & (~x7 ^ ~x8)))) | (~x0 & ((x6 & ~x7 & ~x8) | (x3 & ~x6 & (~x7 ^ x8)))))) | (~x0 & ~x5 & ((~x6 & ~x7 & ~x8) | (x3 & x6 & (~x7 ^ x8)))))) | (~x4 & ((x3 & ((~x6 & x8 & (x0 ? (~x5 ^ x7) : (x5 & ~x7))) | (x7 & ~x8 & ~x0 & x6))) | (x6 & ((x0 & ((~x3 & ~x7) | (~x5 & x7 & ~x8))) | (~x7 & x8 & ~x0 & ~x5))))) | (x6 & x7 & x8 & ~x0 & x3 & x5))) | (~x0 & x3 & x4 & x7 & x8 & ~x5 & ~x6))) | (~x1 & ((~x0 & ((~x3 & ((~x6 & (x2 ? ((~x5 & x7 & x8) | (~x7 & (x8 ? x5 : x4))) : (x4 ? (x7 & ~x8) : (x5 & x8)))) | (x2 & ((~x4 & ~x8 & (x5 ? (x6 & ~x7) : (~x7 | (x6 & x7)))) | (x5 & x6 & x8 & (x7 | (x4 & ~x7))))))) | (x2 & ((~x4 & ((x5 & ~x6 & ~x8 & (x7 | (x3 & ~x7))) | (x3 & x6 & (x7 ? x8 : ~x5)))) | (~x5 & x7 & x8 & x3 & x4))) | (~x2 & ((x4 & ((~x7 & x8 & x5 & x6) | (x3 & (x5 ? (~x6 & ~x8) : (x6 & x8))))) | (x3 & ~x5 & ~x6 & ~x7 & x8))) | (~x6 & x7 & x8 & x3 & x4 & x5))) | (x0 & (x3 ? ((x8 & ((~x2 & ((~x4 & ~x5 & x6) | (~x6 & x7 & x4 & x5))) | (~x7 & (x4 ? (~x5 & ~x6) : x5)))) | (~x6 & x7 & ~x8 & ((~x4 & x5) | (~x2 & x4 & ~x5)))) : ((~x8 & ((~x5 & ((~x6 & ~x7 & x2 & x4) | (x6 & x7 & ~x2 & ~x4))) | (x5 & ((x2 & ~x4 & (~x6 | (x6 & x7))) | (x6 & x7 & ~x2 & x4))) | (x6 & ~x7 & ~x2 & x4))) | (x7 & ((~x2 & ((~x5 & ~x6) | (x4 & x5 & x8))) | (x2 & x4 & ~x5 & ~x6 & x8)))))) | (~x2 & x3 & ~x4 & x7 & ~x8 & ~x5 & ~x6))) | (x2 & x5 & ~x6 & x8 & ((~x0 & x3 & ~x4 & x7) | (x4 & ~x7 & x0 & ~x3)));
  assign z18 = x1 ? (x0 ? ((x6 & (x2 ? (~x3 & ((~x4 & (x7 ? x5 : x8)) | (~x7 & ~x8 & x4 & x5))) : (x3 ? ((x7 & ~x8 & x4 & x5) | (~x7 & x8 & ~x4 & ~x5)) : (~x7 & (x4 ? (~x5 & x8) : (x5 & ~x8)))))) | (x5 & ((~x2 & x3 & x7 & x8 & (~x4 | (x4 & ~x6))) | (x2 & ~x3 & ~x4 & ~x6 & ~x7 & ~x8)))) : (~x3 & ((~x4 & ((~x6 & ((x2 & ~x8 & (~x5 ^ x7)) | (~x7 & x8 & ~x2 & x5))) | (x6 & x7 & ~x8 & ~x2 & ~x5))) | (x2 & x4 & ~x7 & x8 & (~x5 ^ ~x6))))) : ((~x4 & ((x6 & ((~x2 & ((~x0 & x5 & ~x8 & (x3 ^ x7)) | (x7 & x8 & x0 & x3))) | (x0 & x2 & ~x5 & (x3 ? (x7 & x8) : (~x7 & ~x8))))) | (~x7 & x8 & ~x5 & ~x6 & ~x0 & x2 & x3))) | (x2 & ((x0 & ~x8 & ((x3 & x4 & (x5 ? (~x6 & x7) : (x6 & ~x7))) | (~x3 & ~x5 & ~x6 & x7))) | (x5 & ~x6 & ~x7 & ~x0 & ~x3 & x4))));
  assign z19 = (~x0 & ((~x2 & (((~x6 ^ x7) & ((x5 & x8 & ~x1 & ~x4) | (x1 & ~x3 & x4 & ~x5 & ~x8))) | (x1 & ((~x7 & (x3 ? ((x5 & x6 & x8) | (~x4 & ~x5 & ~x6)) : ((x4 & x6 & x8) | (~x8 & (x5 ? ~x6 : ~x4))))) | (x4 & ((~x3 & x5 & x7 & (x6 ^ ~x8)) | (~x6 & x8 & x3 & ~x5))))) | (~x3 & ~x7 & ((~x1 & x4 & ~x5) | (x6 & ~x8 & ~x4 & x5))) | (~x1 & x3 & ((~x4 & (x5 ? (~x8 & (~x6 | (x6 & x7))) : (x6 & x7))) | (~x6 & x7 & ~x8 & x4 & ~x5))))) | (x2 & (x3 ? ((x8 & ((x1 & ((x5 & x6 & x7) | (~x6 & ~x7 & ~x4 & ~x5))) | (~x6 & x7 & ~x1 & ~x4))) | (~x1 & ~x4 & ~x8 & (x5 ? (~x6 & ~x7) : (x6 & x7)))) : (x6 ? ((x8 & ((x4 & ~x5 & x7) | (~x1 & (x7 ? ~x4 : x5)))) | (x1 & ~x4 & (x5 ? (~x7 | (x7 & ~x8)) : ~x8))) : ((x1 & (x4 ? (x8 & (~x5 ^ x7)) : (x5 & x7))) | (x7 & ~x8 & ~x1 & ~x5) | (~x4 & (x5 ? ~x7 : x8)))))) | (x7 & ~x8 & ((~x1 & ~x3 & x4 & ~x5 & x6) | (x1 & x3 & ~x4 & x5 & ~x6))))) | (x0 & ((~x2 & (x1 ? (x5 ? ((~x4 & (x8 ? ~x3 : x7)) | (~x6 & ~x8 & x3 & x4)) : (x3 ? ((x4 & ~x8 & (x7 | (x6 & ~x7))) | (x7 & x8 & ~x4 & ~x6)) : (x4 ? (~x6 & x7) : (x6 & ~x7)))) : ((x8 & (x3 ? ((~x4 & ~x6 & x7) | (x6 & ~x7 & x4 & ~x5)) : (x5 & (x7 ? x6 : ~x4)))) | (~x6 & x7 & ~x8 & ~x4 & x5) | (~x3 & ((~x6 & ~x7 & ~x4 & ~x5) | (x4 & ((~x5 & x6 & x7) | (~x6 & ~x7 & ~x8)))))))) | (x2 & ((~x1 & (x5 ? ((~x4 & (x3 ? (x6 ? ~x8 : (x7 & x8)) : (x7 & ~x8))) | (~x3 & x4 & (x6 ? x8 : x7))) : (x3 ? (~x4 & (x6 ? (~x7 & x8) : (x8 | (x7 & ~x8)))) : ((x6 & ~x7) | (x4 & ~x6 & ~x8))))) | (~x3 & ((x1 & (x4 ? ((~x7 & x8 & ~x5 & x6) | (x7 & ~x8 & x5 & ~x6)) : ((x7 & ~x8 & ~x5 & x6) | (~x7 & (x5 ? (x6 ^ x8) : ~x8))))) | (x7 & x8 & x4 & ~x5))))) | (~x1 & ~x4 & ~x7 & ((x3 & (x5 ? (x6 & x8) : (~x6 & ~x8))) | (x6 & ~x8 & ~x3 & x5))))) | (~x3 & x7 & ((~x1 & x4 & ((~x6 & x8 & ~x2 & ~x5) | (x6 & ~x8 & x2 & x5))) | (~x5 & x6 & x8 & x1 & x2 & ~x4))) | (~x7 & x8 & x5 & ~x6 & x3 & x4 & ~x1 & ~x2);
  assign z20 = (x8 & (x4 ? ((~x0 & (x3 ? (x7 & ((x2 & (~x5 | (x5 & ~x6))) | (x5 & x6 & ~x1 & ~x2))) : ((x1 & ((x6 & x7 & x2 & x5) | (~x2 & ~x6 & ~x7))) | (x2 & ((~x5 & x6 & ~x7) | (~x1 & x5 & x7)))))) | (x0 & ((x5 & ~x6 & ~x2 & ~x3) | (x1 & (x2 ? (~x3 & ~x7 & (~x6 | (x5 & x6))) : (x5 & x6))))) | (~x1 & ~x2 & ~x3 & x5 & x6 & ~x7)) : (x6 ? (x0 ? ((~x1 & ((x2 & x5 & x7) | (~x2 & x3 & ~x5 & ~x7))) | (~x5 & x7 & ~x2 & ~x3)) : (x2 & (x1 ? (~x5 & ~x7) : (x3 ? x7 : (x5 & ~x7))))) : ((x1 & ((~x0 & x3 & (x7 ? ~x2 : x5)) | (x0 & ~x2 & ~x3 & ~x5 & ~x7))) | (x0 & ((~x1 & x5 & ~x7 & (x3 | (x2 & ~x3))) | (~x5 & x7 & x2 & ~x3))))))) | (~x8 & ((x4 & ((~x3 & (x6 ? ((x1 & ((x5 & x7 & x0 & x2) | (~x5 & ~x7 & ~x0 & ~x2))) | (x0 & ~x1 & x7 & (x2 ^ x5))) : ((~x0 & (x1 ? (x2 & x7) : (~x5 & ~x7))) | (~x5 & ~x7 & x0 & x1)))) | (~x2 & ((x3 & (x0 ? (~x1 & ((x6 & ~x7) | (x5 & ~x6 & x7))) : (x1 & ~x7 & (~x6 | (x5 & x6))))) | (~x1 & ~x6 & x7 & (x0 ^ x5)))) | (x0 & ~x1 & x2 & ~x7 & ((x5 & x6) | (x3 & ~x5 & ~x6))))) | (~x4 & ((x7 & (x3 ? ((~x0 & x2 & (x1 ? (x5 ^ ~x6) : (x5 & ~x6))) | (~x2 & ~x5 & ~x6)) : (x0 ? ((~x1 & ~x2 & ~x5) | (x5 & ~x6 & x1 & x2)) : ((~x1 & x2 & x6) | (~x5 & ~x6 & x1 & ~x2))))) | (~x0 & ~x1 & x2 & ~x5 & ~x7 & (~x6 | (x3 & x6))))) | (~x0 & x1 & ~x2 & x6 & x7 & x3 & ~x5))) | (~x0 & ~x1 & ~x2 & x3 & ~x5 & ~x7 & (~x4 ^ x6));
  assign z21 = x8 ? (x3 ? (x1 ? ((~x4 & ((x2 & ((x0 & (x5 ? (~x6 & ~x7) : x7)) | (~x6 & x7 & ~x0 & x5))) | (~x5 & x6 & ~x7 & ~x0 & ~x2))) | (x5 & ~x6 & ~x7 & ~x0 & ~x2 & x4)) : ((~x0 & ((~x2 & x4 & x5 & ~x6 & x7) | (~x5 & x6 & ~x7 & x2 & ~x4))) | (~x2 & x4 & x5 & x6 & ~x7))) : (x0 ? (~x6 & ((~x1 & ~x5 & (x2 ? (x4 & ~x7) : (~x4 & x7))) | (x1 & x2 & x4 & x5 & x7))) : ((x4 & ~x5 & ~x6 & ~x1 & x2) | (x5 & x6 & x7 & ~x2 & ~x4)))) : ((x1 & (x0 ? (x2 & ~x7 & ((x3 & ~x5 & (~x4 | (x4 & x6))) | (x5 & ~x6 & ~x3 & ~x4))) : ((x4 & (x2 ? (~x7 & (x3 | (~x3 & x6))) : ((~x3 & x5 & x6) | (~x6 & x7 & x3 & ~x5)))) | (~x5 & x6 & x7 & x2 & x3 & ~x4)))) | (x0 & ((x2 & x3 & ~x6 & (x4 ? (~x5 & ~x7) : (x5 & x7))) | (x4 & x6 & ~x7 & ~x1 & ~x2 & ~x3))));
  assign z22 = (x0 & ((x5 & ((~x8 & ((x1 & ((x6 & (x2 ? (~x3 & x4) : (x7 & (x3 ^ ~x4)))) | (x2 & ~x4 & (x7 ? ~x6 : x3)) | (~x2 & x3 & x4 & ~x6 & ~x7))) | (~x1 & ((x7 & (x2 ? (x3 ? x6 : ~x4) : (~x4 ^ x6))) | (x6 & ~x7 & (~x3 | (x3 & x4))))) | (x2 & ~x3 & x4 & ~x6 & x7))) | (x8 & ((x1 & ((x7 & (x2 ? (x3 ? (~x4 & ~x6) : x6) : (x3 & x4))) | (~x3 & ((~x2 & (x6 ? x4 : ~x7)) | (~x6 & ~x7 & x2 & ~x4))))) | (~x4 & ((~x2 & x3 & x7) | (~x1 & ~x7 & (x2 ? (x3 & x6) : ~x3)))) | (~x1 & ((~x3 & ((x6 & x7) | (x2 & x4 & (~x6 | (x6 & ~x7))))) | (~x6 & x7 & ~x2 & x4))))) | (~x1 & ~x6 & ((~x4 & (x2 ? (~x3 ^ x7) : (x3 & ~x7))) | (~x2 & ~x3 & x4 & ~x7))))) | (~x5 & (x1 ? (x2 ? (x3 ? (~x7 & (x4 ? (x6 & ~x8) : x8)) : (x4 & x8)) : ((x6 & ((~x4 & ~x7 & ~x8) | (x3 & (x4 ^ x8)))) | (~x6 & x7 & ~x8) | (~x3 & ~x7 & (x4 ? (~x6 & ~x8) : x8)))) : ((~x2 & ((~x8 & ((x3 & (x4 ? x7 : ~x6)) | (x4 & x6 & ~x7) | (~x3 & (~x6 | (x6 & x7))))) | (~x4 & x7 & x8) | (x4 & ((x6 & x7 & x8) | (x3 & ~x6 & ~x7))))) | (x2 & ((~x4 & ((~x6 & x7) | (x3 & (x6 ? x8 : ~x7)))) | (~x3 & ((x6 & ~x7) | (x4 & (x7 ? x8 : ~x6)))))) | (x3 & x4 & x6 & ~x7 & x8)))) | (~x3 & ((x2 & ~x8 & ((x6 & x7 & ~x1 & x4) | (~x6 & ~x7 & x1 & ~x4))) | (x1 & ~x2 & x7 & x8 & (~x4 ^ ~x6)))) | (~x1 & ~x2 & x3 & ~x4 & x6 & (~x7 ^ ~x8)))) | (~x0 & ((~x3 & ((x4 & ((~x1 & (x2 ? (x7 ? x8 : (~x6 | (x5 & x6))) : ((x7 & ~x8) | (~x5 & ~x6 & x8)))) | (x1 & ((x2 & (x6 ? (~x7 ^ x8) : (x5 ? (x7 & x8) : (~x7 | (x7 & ~x8))))) | (x5 & ~x6 & (x7 ? ~x8 : ~x2)))) | (x6 & x7 & ~x8 & x2 & ~x5))) | (x2 & ((~x4 & ((x1 & (~x6 | (x5 & x6 & ~x7))) | (x5 & ~x8 & (x7 ? x6 : ~x1)) | (~x1 & x8 & (x6 ? x7 : ~x5)))) | (~x6 & x7 & ~x8 & ~x1 & ~x5))) | (~x4 & ((x5 & ((~x1 & ((~x6 & ~x7 & x8) | (~x2 & x6 & ~x8))) | (~x7 & x8 & x1 & ~x2))) | (x1 & ~x5 & ((x6 & ~x7) | (~x2 & (x8 ? ~x6 : x7)))))) | (x1 & ~x2 & x5 & x6 & (~x7 ^ x8)))) | (x3 & ((~x4 & (x6 ? ((x1 & ((~x2 & ((~x7 & x8) | (~x5 & x7 & ~x8))) | (x7 & ~x8 & x2 & x5))) | (~x1 & ((~x2 & ~x7 & ~x8) | (x5 & x8 & (~x7 | (x2 & x7))))) | (x2 & ~x5 & (~x7 ^ ~x8))) : ((x1 & (x2 ? (x5 & x8) : ~x5)) | (~x1 & ~x5 & ~x7) | (x7 & ~x8 & x2 & x5)))) | (x4 & (x7 ? ((x8 & (x6 ? (x1 ? (~x5 | (x2 & x5)) : (~x2 & x5)) : (x2 ? x5 : ~x1))) | (x6 & ~x8 & ~x2 & ~x5)) : ((x1 & (x2 ? ~x8 : (x5 & x6))) | (~x2 & x5 & ~x6)))) | (~x1 & x7 & (x2 ? (~x5 & x8) : (~x8 & (x5 ^ ~x6)))))) | (~x2 & ((x4 & ~x5 & (x1 ? (~x6 | (x6 & ~x7 & x8)) : (x6 & ~x7))) | (x6 & x7 & x8 & ~x1 & ~x4 & x5))))) | (x7 & ((x4 & ((x1 & ~x5 & ((~x6 & x8 & x2 & x3) | (x6 & ~x8 & ~x2 & ~x3))) | (~x2 & x3 & x5 & ~x6 & ~x8))) | (x1 & x2 & ~x4 & ~x5 & (x3 ? (~x6 & ~x8) : x6)))) | (~x7 & x8 & x5 & x6 & ~x1 & ~x2 & x4);
  assign z23 = (~x7 & ((x0 & ((x1 & (x2 ? ((~x4 & ((~x6 & x8 & ~x3 & ~x5) | (x3 & (x5 ? x8 : (x6 & ~x8))))) | (~x3 & x4 & x5 & x6 & x8)) : (~x8 & ((x3 & (x4 ? (~x5 & ~x6) : x5)) | (~x3 & x4 & x5) | (~x4 & ~x5 & ~x6))))) | (~x1 & (x8 ? ((~x5 & ((~x2 & (x3 ? (~x4 & ~x6) : (x4 & x6))) | (x4 & ~x6 & x2 & x3))) | (x2 & x5 & x6 & (x3 ^ ~x4))) : ((~x2 & ~x3 & ~x4 & ~x5 & x6) | (x2 & x3 & x4 & x5 & ~x6)))) | (x5 & ~x6 & ~x8 & ~x2 & ~x3 & ~x4))) | (~x0 & ((~x1 & ((x2 & ((x3 & x5 & ~x6) | (x6 & ~x8 & ~x3 & ~x5))) | (~x2 & ((~x3 & (x4 ? (x5 & ~x8) : ~x5)) | (~x5 & x6 & x3 & ~x4))) | (x3 & x4 & ~x8 & (x5 ^ ~x6)))) | (x4 & ((x1 & ((x2 & x8 & (x3 ? (x5 & ~x6) : x6)) | (~x2 & ~x3 & ~x5 & x6 & ~x8))) | (x2 & x3 & x8 & (~x5 | (x5 & x6))))) | (x6 & ~x8 & ~x4 & x5 & x1 & x2 & x3))) | (x1 & x2 & x3 & ~x6 & ~x8 & ~x4 & ~x5))) | (x7 & ((~x0 & ((~x2 & (x4 ? (x8 & ((~x1 & x6 & (~x3 | (x3 & ~x5))) | (~x3 & x5 & ~x6))) : ((x1 & ((~x5 & x6 & x8) | (~x3 & x5 & ~x8))) | (~x1 & x3 & ~x5 & ~x6 & x8)))) | (~x1 & x2 & ((x3 & (x5 ? (x4 ? ~x8 : (~x6 & x8)) : (~x6 & ~x8))) | (~x6 & ~x8 & ~x3 & x5))))) | (x0 & (x1 ? (x6 & ((x3 & ~x4 & (x5 ? x2 : ~x8)) | (~x2 & ~x3 & x4 & ~x5 & x8))) : ((~x2 & ((x3 & x4 & ~x5 & ~x6 & x8) | (~x3 & ~x4 & x5 & x6 & ~x8))) | (x4 & ((x2 & ~x5 & (x6 ? x3 : ~x8)) | (x3 & x5 & x6 & x8))) | (x2 & ~x3 & ~x4 & ~x5 & x6 & ~x8)))) | (x1 & x2 & x3 & ~x4 & ~x5 & x8))) | (~x0 & ~x1 & x2 & x3 & x6 & ~x8 & (~x4 ^ ~x5));
  assign z24 = x0 ? (~x5 & ((x2 & (x7 ? ((~x8 & ((x1 & ~x6 & (x3 ^ ~x4)) | (x4 & x6 & ~x1 & x3))) | (~x1 & ~x3 & ~x4 & x6 & x8)) : ((x1 & x4 & (x8 ? x3 : ~x6)) | (~x1 & ~x3 & ~x4 & ~x6 & ~x8)))) | (x7 & x8 & x4 & x6 & x1 & ~x2 & ~x3))) : (x1 ? (~x2 & x3 & ((x7 & ~x8 & x5 & x6) | (x4 & ((x7 & x8 & x5 & ~x6) | (~x7 & ~x8 & ~x5 & x6))))) : ((x7 & (x2 ? (x3 & x5 & (x6 ? ~x8 : (x4 ^ x8))) : (~x3 & ((~x4 & ~x5) | (x6 & x8 & x4 & x5))))) | (~x8 & ((x2 & x3 & ((x5 & ~x6 & ~x7) | (x4 & (~x5 | (x5 & x6 & ~x7))))) | (~x2 & ~x3 & x4 & x5 & ~x7)))));
  assign z25 = (x0 & (x1 ? (x2 ? (x3 & ((~x4 & ((x7 & x8 & ~x5 & ~x6) | ((~x6 ^ x7) & (x5 ^ ~x8)))) | (x6 & ~x7 & ~x8 & x4 & ~x5))) : ((x6 & x7 & x8 & ~x3 & x4 & ~x5) | (x3 & ~x4 & x5 & ~x6 & ~x7 & ~x8))) : (x3 & x4 & ((x6 & ((x5 & x7 & x8) | (x2 & (x5 ? (~x7 & x8) : (x7 & ~x8))))) | (x2 & ~x5 & ~x6 & ~x7 & x8))))) | (x7 & x8 & x4 & ~x5 & ~x0 & ~x1 & ~x2 & x3);
  assign z26 = x1 ? (~x5 & ((~x6 & ((~x4 & (x0 ? (~x3 & (x2 ? (~x7 & x8) : ~x8)) : (x2 & x3 & (~x7 ^ x8)))) | (x4 & ~x7 & ~x8 & x0 & ~x2 & ~x3))) | (~x0 & x2 & ~x3 & ~x7 & x8 & x4 & x6))) : (x4 ? (~x5 & ((x2 & ((x0 & ~x6 & ~x8 & (~x3 ^ x7)) | (x6 & x7 & x8 & ~x0 & ~x3))) | (~x0 & ~x2 & x3 & ~x7 & ~x8))) : (x0 ? (~x3 & ~x8 & ((x6 & x7 & x2 & ~x5) | (~x6 & ~x7 & ~x2 & x5))) : (x3 & x8 & ((x6 & x7 & ~x2 & x5) | (~x6 & ~x7 & x2 & ~x5)))));
  assign z27 = (~x0 & ((x5 & ((~x1 & ((x4 & ((~x8 & (x2 ? (x7 ? x3 : x6) : (~x6 & x7))) | (~x6 & ~x7) | (x8 & ((x3 & (~x6 ^ ~x7)) | (~x2 & x6 & x7))))) | (x2 & ((~x3 & (x7 ? x8 : ~x4)) | (x7 & x8 & x3 & x6))) | (x3 & ~x4 & (~x6 | (x6 & x7 & ~x8))))) | (x1 & ((~x7 & ((~x2 & ~x3 & ~x6) | (x3 & x4 & x6))) | (x7 & ((x6 & ((x4 & ~x8) | (x3 & (x2 ? (x4 ^ ~x8) : x8)))) | (~x2 & ~x3 & ~x4 & x8))) | (x3 & ~x6) | (x2 & ((~x3 & ~x6) | (x6 & x8 & x3 & ~x4))))) | (x3 & ~x4 & x6 & ~x7 & (~x2 | (x2 & ~x8))))) | (~x5 & ((x6 & ((x2 & ((~x8 & (x1 ? (x3 ? ~x7 : x4) : (x3 & x7))) | (x7 & x8 & x3 & x4) | (~x1 & (x3 ? (x4 & ~x7) : (~x4 & x8))))) | (x1 & ((x3 & ((x4 & x7 & ~x8) | (~x2 & ~x7))) | (~x2 & x7 & (x8 ? x4 : ~x3)))))) | (~x6 & ((x1 & ~x2 & (~x4 | (x3 & x4))) | (~x1 & ~x3 & x4) | (x2 & (x3 ^ ~x4)))) | (x3 & ((x2 & ~x4 & (x1 ? (x7 & ~x8) : (~x7 ^ x8))) | (~x1 & ~x2 & x4 & ~x7 & x8))))) | (x6 & ((~x4 & ((x2 & (x1 ? ~x3 : (x3 ? (~x7 & x8) : (x7 & ~x8)))) | (x1 & ~x2 & (x3 ? (x7 & ~x8) : ~x7)))) | (~x3 & x4 & ((~x1 & ((x7 & ~x8) | (x2 & ~x7 & x8))) | (~x2 & ~x7) | (x7 & x8 & x1 & x2))))) | (~x2 & ~x3 & ((~x1 & ~x4) | (~x6 & x7 & ~x8 & x1 & x4))))) | (x0 & ((x1 & ((~x5 & (x2 ? ((x6 & ((~x3 & x4) | (x7 & x8 & x3 & ~x4))) | (~x6 & (x3 ? (x4 & (~x7 ^ x8)) : (~x4 & ~x8))) | (x7 & x8 & ~x3 & ~x4)) : (x4 ? ((x6 & ~x7) | (x3 & (x8 ? ~x6 : x7))) : (x3 ? (~x6 | (x6 & ~x7)) : (x6 | (~x6 & x8)))))) | (x3 & ((x5 & ((~x4 & (x2 ? (x6 ? (~x7 & x8) : (~x7 ^ x8)) : (x8 ? ~x6 : x7))) | (~x2 & (x6 ? ((~x7 & x8) | (x4 & (~x8 | (x7 & x8)))) : x4)))) | (~x4 & ((x2 & ~x8 & (~x6 ^ ~x7)) | (x7 & x8 & ~x2 & x6))))) | (~x3 & ((x4 & ((x6 & x7 & x2 & x5) | (~x2 & ((x7 & ~x8) | (x5 & ~x6 & x8))))) | (x2 & ~x4 & (x6 ? (~x7 | (x7 & ~x8)) : x5)))))) | (~x3 & ((~x1 & (x2 ? ((~x4 & (~x6 | (x5 & x6 & ~x8))) | (x7 & ((x6 & x8) | (x4 & ~x5 & ~x8))) | (~x5 & x6 & ~x7) | (x4 & (x5 ? (x6 & ~x7) : (~x6 & x8)))) : ~x5)) | (x5 & (x2 ? (x4 & ~x6) : ((x6 & (~x7 | (x7 & x8))) | (~x4 & (x8 ? ~x6 : x7))))))) | (~x1 & ((x3 & (x4 ? ((~x7 & (((~x5 | (x5 & x6)) & (~x2 | (x2 & ~x8))) | (x2 & x5 & ~x6))) | (x2 & ~x6 & x7 & (x8 | (x5 & ~x8)))) : (x5 | (x2 & ~x5)))) | (x4 & x5 & (x6 ? (x7 & ~x8) : ~x2)))) | (x3 & x4 & ~x5 & x6 & x8 & (~x2 ^ ~x7)))) | (~x5 & ((~x2 & ((~x1 & x3 & (~x4 | (x4 & x7 & ~x8))) | (x1 & ~x3 & x4 & ~x6 & x8))) | (x1 & x2 & ((~x3 & x4 & ~x6) | (~x7 & x8 & x3 & ~x4))))) | (x1 & x2 & ~x3 & x6 & ~x7 & x4 & x5);
  assign z28 = x1 ? (x0 ? ((x3 & ~x8 & (((x4 ? (~x5 & ~x6) : (x5 & x6)) & (x2 ^ ~x7)) | (~x2 & ~x4 & ~x5 & x6 & x7))) | (x2 & ~x3 & ~x4 & x7 & x8 & x5 & x6)) : (~x2 & x7 & ((~x3 & x5 & (x4 ? (~x6 & x8) : ~x8)) | (x6 & x8 & ~x4 & ~x5)))) : ((x2 & ((~x3 & ((~x0 & ~x8 & ((x5 & ~x6 & x7) | (x6 & ~x7 & ~x4 & ~x5))) | (x6 & ~x7 & x8 & x0 & ~x4 & x5))) | (~x0 & x3 & ~x4 & x7 & ~x8 & ~x5 & ~x6))) | (x7 & x8 & ~x5 & x6 & ~x3 & x4 & ~x0 & ~x2));
  assign z29 = (x0 & ((x3 & ((x4 & ((x1 & ((~x6 & (((~x7 | (x7 & x8)) & (x2 ^ x5)) | (~x2 & ~x5 & x8))) | (~x2 & x6 & ((x7 & x8) | (x5 & ~x7 & ~x8))))) | (~x5 & ((~x2 & (x6 ? (x7 & ~x8) : ~x1)) | (~x1 & x2 & (x7 ? x8 : (~x8 | (x6 & x8)))))) | (~x1 & x5 & ~x6 & ((x7 & ~x8) | (x2 & (~x7 | (x7 & x8))))))) | (~x4 & ((x1 & (x6 ? (x2 ? ((~x7 & ~x8) | (~x5 & x7 & x8)) : (x5 ? (x7 & ~x8) : ~x7)) : (x2 ? ((x7 & ~x8) | (x5 & (~x7 ^ x8))) : (x5 & x8)))) | (~x5 & (x2 ? ~x1 : (~x6 & x8))) | (x7 & x8 & ~x2 & x6) | (~x1 & ((~x2 & x7 & ~x8) | (x5 & ((~x6 & ~x7) | (x2 & (~x6 ^ ~x7)))))))) | (~x2 & (x1 ? ((~x6 & x7 & ~x8) | (~x7 & x8 & x5 & x6)) : (x6 & ~x7))))) | (x6 & (((x2 ? (~x3 & ~x4) : (x4 & ~x5)) & (x1 ? ~x7 : (x7 & x8))) | (~x3 & (x1 ? (x2 ? (x4 ? (~x5 | (x5 & (~x8 | (x7 & x8)))) : (x7 & ~x8)) : (~x4 | (x4 & x5 & x8))) : (x2 ? ((x4 & (x7 | (x5 & ~x7))) | (~x5 & ~x7) | (~x4 & x5 & ~x8)) : ((~x4 & (x8 ? ~x5 : x7)) | (x5 & (~x7 | (x7 & x8))) | (x4 & ~x5 & ~x8))))) | (~x2 & x4 & x5 & x7 & ~x8))) | (~x6 & (x1 ? (~x3 & (x2 ? (x4 ? (x5 & ~x7) : (x5 | (~x5 & ~x8))) : (x5 | (~x5 & x8)))) : ((~x3 & (x2 ? (~x4 | (x4 & (x5 | (~x5 & x8)))) : (~x5 | (x5 & (x8 ? ~x4 : x7))))) | (~x2 & x4 & x5 & (~x7 | (x7 & x8)))))) | (x1 & ~x3 & ~x5 & x7 & (x2 ? (~x4 & x8) : (x4 & ~x8))))) | (~x0 & ((~x3 & ((x1 & ((x2 & (~x4 | (x4 & x6 & ~x8))) | (x7 & x8 & x4 & x6) | (~x2 & ((x5 & ((~x6 & ~x7) | (~x4 & x7 & x8))) | (x6 & ~x7) | (~x5 & (~x6 | (x6 & x7 & ~x8))))))) | (~x1 & ((~x2 & (~x4 | (x4 & ~x6))) | (x6 & ((x4 & (~x7 | (x7 & ~x8))) | (x2 & ~x4 & (x8 ? ~x5 : x7)))) | (x2 & (x5 ? (x7 ? x8 : ~x4) : ~x6)))) | (x5 & ~x6 & ~x7 & x2 & x4))) | (x3 & ((~x2 & (((x1 ? ~x4 : x5) & (~x6 | (x6 & (~x7 | (x7 & ~x8))))) | (x1 & ((x7 & x8 & x5 & x6) | (x4 & (~x5 | (x5 & ~x7))))) | (~x1 & ~x5 & (x7 ? ~x8 : (~x4 | (x4 & x8)))))) | (x2 & ((~x8 & ((~x5 & (x1 ? ((~x4 & x7) | (x6 & (~x7 | (x4 & x7)))) : (x4 | (~x4 & ~x7)))) | (~x1 & x5 & ~x6) | (x1 & ((x5 & x6 & x7) | (x4 & (~x6 | (x5 & x6 & ~x7))))))) | (x8 & (x4 ? (x7 & (~x5 | (x5 & (~x6 | (x1 & x6))))) : ((~x1 & ~x6 & x7) | (x6 & (x1 ? (x7 | (x5 & ~x7)) : ~x7))))) | (x5 & ~x6 & x1 & ~x4))) | (~x1 & x6 & x7 & x8 & (~x4 ^ x5)))) | (x5 & x7 & ~x8 & x1 & ~x2 & x4))) | (x2 & ((x3 & (x1 ? (~x5 & ~x7 & x8 & (~x4 | (x4 & x6))) : (x5 & x6 & (x4 ? ~x8 : x7)))) | (x1 & ~x3 & x4 & ~x6 & (~x5 | (x5 & x7)))));
  assign z30 = (~x3 & ((~x6 & (x2 ? ((x7 & ((x8 & ((x5 & (x0 ? (~x1 | (x1 & x4)) : ~x4)) | (x1 & x4 & ~x5))) | (~x0 & ~x1 & ~x5 & ~x8))) | (x1 & (x4 ? (x5 & ~x7) : (x0 ? (x5 ? x8 : (~x7 & ~x8)) : (~x5 & x8)))) | (~x0 & ~x4 & x5 & ~x7 & ~x8)) : ((~x0 & ((~x7 & ((x1 & ~x8 & (~x4 | (x4 & ~x5))) | (~x1 & x4 & x5 & x8))) | (x5 & ~x8 & ~x1 & ~x4))) | (x0 & ((~x1 & ((~x5 & ~x7) | (~x4 & x5 & x8))) | (x7 & ((x5 & ~x8) | (x1 & ~x4 & x8))))) | (~x1 & x4 & ~x5 & x7 & x8)))) | ((x0 ? (x2 & ~x5) : (x5 & x6)) & ((~x7 & x8 & ~x1 & ~x4) | (x7 & ~x8 & x1 & x4))) | (~x5 & ((x8 & ((x6 & ((x4 & ((~x0 & x1 & ~x2) | (x7 & (x0 ? (~x1 | (x1 & x2)) : x2)))) | (~x0 & ~x1 & x2 & ~x7))) | (x0 & x1 & x2 & ~x4 & x7))) | (x4 & ((~x0 & ~x2 & ((x6 & x7 & ~x8) | (~x1 & ~x7))) | (x6 & ~x7 & x0 & x2))))) | (x0 & ((x5 & ((x6 & ((x7 & ((~x2 & ~x4 & x8) | (x1 & ~x8 & (x2 ^ x4)))) | (x4 & x8 & ~x1 & x2))) | (x4 & x7 & ~x8 & ~x1 & x2))) | (~x2 & ~x4 & x6 & ((~x7 & x8) | (x1 & x7 & ~x8))))) | (~x0 & x1 & x2 & ~x4 & ((x5 & ~x7 & x8) | (x6 & (~x8 | (x7 & x8))))))) | (x3 & ((x7 & (x2 ? ((x4 & ((~x1 & ((x0 & ~x6 & (x8 | (x5 & ~x8))) | (x6 & x8 & ~x0 & x5))) | (~x0 & x1 & ~x8))) | (~x1 & ~x4 & ((~x5 & ~x6 & x8) | (x0 & (x5 ? (x6 & x8) : ~x8))))) : ((~x4 & ((x0 & ((~x1 & ~x6 & x8) | (x6 & ~x8 & x1 & x5))) | (~x0 & ((x5 & x6 & x8) | (~x1 & (x5 ? ~x8 : x6)))) | (~x6 & ~x8 & x1 & x5))) | (x1 & x4 & ((x5 & (x0 ? (~x6 & ~x8) : (x6 & x8))) | (x0 & ~x5 & (~x8 | (x6 & x8)))))))) | (~x7 & (x4 ? ((x0 & ((~x1 & x2 & (x5 ? (~x6 & x8) : ~x8)) | (~x2 & x5 & (~x6 | (x1 & x6))))) | (~x5 & ~x6 & x8 & ~x0 & ~x1 & ~x2)) : (x5 ? ((~x0 & ((~x2 & ~x6) | (x1 & ~x8 & (~x2 ^ ~x6)))) | (x0 & x1 & ~x2 & x8)) : (x0 ? (~x1 & (x2 | (~x2 & ~x8))) : (x1 & (x2 ? (x6 ^ x8) : ~x8)))))) | (~x4 & ((x2 & ((~x1 & ((x0 & x5 & (x6 ^ x8)) | (x6 & ~x8 & ~x0 & ~x5))) | (~x0 & x1 & x5 & x6 & x8))) | (x0 & x1 & ~x2 & ~x5 & ~x6 & x8))))) | (~x2 & ((x5 & ((~x0 & x8 & ((~x4 & ~x6 & x7) | (x6 & ~x7 & x1 & x4))) | (x6 & ~x7 & ~x8 & x0 & ~x1 & ~x4))) | (x0 & x1 & x4 & ~x5 & (x6 ? ~x7 : x8))));
  assign z31 = (x2 & ((~x1 & ((~x5 & ((~x3 & ((~x0 & ((x6 & ~x7 & x8) | (~x4 & ~x6 & ~x8))) | (x7 & ~x8 & x4 & ~x6) | (~x7 & x8 & x0 & ~x4))) | (x0 & x3 & (x4 ? ((x6 & (~x7 ^ x8)) | (x7 & ~x8) | (~x6 & ~x7)) : (~x6 ^ ~x7))) | (x6 & x7 & ~x8 & ~x0 & ~x4))) | (x6 & x7 & x8 & x3 & x4 & x5) | (x0 & ((x4 & ((x7 & x8 & ~x3 & x6) | (x5 & ((x3 & ((~x7 & x8) | (~x6 & x7 & ~x8))) | (x7 & ~x8 & ~x3 & x6) | (~x6 & (~x7 ^ x8)))))) | (x3 & ~x4 & ((x6 & ~x8 & (x7 | (x5 & ~x7))) | (x5 & (x7 ? x8 : ~x6)))) | (x6 & ~x7 & x8 & ~x3 & x5))))) | (x1 & ((~x0 & (x3 ? (x4 ? ((x7 & ~x8) | (~x6 & ~x7 & x8)) : (x5 ? (x6 ? x8 : (~x7 & ~x8)) : (~x6 & ~x7))) : (~x4 & ((x6 & (~x8 | (x7 & x8))) | (x8 & (x5 ? ~x7 : ~x6)))))) | (x0 & (x5 ? ((~x4 & ((x8 & (x3 ? (~x7 | (x6 & x7)) : ~x6)) | (x6 & (x7 ? ~x8 : ~x3)))) | (~x3 & x4 & x8 & (~x6 ^ ~x7))) : ((~x3 & x4 & x7) | (~x4 & ((x3 & ~x8 & (~x7 | (x6 & x7))) | (x7 & x8) | (~x3 & ~x7)))))) | (~x3 & x4 & x5 & ~x6 & ~x7))) | (~x0 & ((~x4 & (x3 ? (~x5 & (x6 ? (~x7 & ~x8) : (x7 & x8))) : (x5 & ~x6 & (~x7 ^ x8)))) | (~x3 & x4 & x6 & x7 & (~x5 ^ ~x8)))) | (~x5 & x6 & ~x7 & x0 & ~x3 & x4))) | (x0 & (x1 ? (~x2 & ((x5 & ((~x4 & ((x3 & ~x7 & ~x8) | (x7 & x8 & ~x3 & x6))) | (~x8 & ((x4 & ~x6 & ~x7) | ((~x3 | (x3 & x4)) & (~x6 ^ ~x7)))) | (x3 & ~x7 & x8 & (x6 | (x4 & ~x6))))) | (~x5 & (((~x7 | (x7 & x8)) & (x6 ? x4 : x3)) | (x4 & (x3 ? (x7 & ~x8) : (~x6 & x8))))) | (~x4 & ((x6 & ((x7 & ~x8) | (~x3 & ~x7 & x8))) | (~x3 & ~x6 & (~x7 ^ x8)))))) : ((~x8 & ((~x3 & x4 & x5 & ~x6 & x7) | (~x2 & x3 & ~x4 & x6 & ~x7))) | (~x2 & (x4 ? (x3 ? (x5 & (x6 ? (x7 & x8) : ~x7)) : (~x5 & (x6 ? x8 : ~x7))) : ((~x3 & (x5 | (~x5 & ~x7))) | (x7 & x8 & x3 & ~x6)))) | (x3 & ~x5 & ~x6 & (x4 ? (x7 & x8) : ~x7))))) | (~x2 & ((~x0 & (x4 ? ((x8 & ((x6 & ((x1 & (x3 ? (x5 & x7) : ~x5)) | (x5 & x7 & ~x1 & ~x3))) | (~x1 & ~x6 & ~x7 & (~x3 ^ ~x5)))) | (~x3 & ((x7 & ~x8 & ~x5 & x6) | (~x7 & ((~x1 & (~x5 | (x5 & x6 & ~x8))) | (~x6 & ~x8 & x1 & ~x5)))))) : ((~x1 & ((~x6 & ~x8 & ~x3 & x5) | (x3 & ((x5 & ~x6 & ~x7) | (x7 & (x5 ? (~x8 | (x6 & x8)) : x6)))))) | (~x6 & ((x5 & x7 & x8) | (x1 & ~x7 & ~x8)))))) | (x1 & x5 & ((x3 & ~x4 & ~x6 & (~x7 ^ ~x8)) | (x6 & x7 & ~x8 & ~x3 & x4))) | (~x1 & ~x3 & x4 & x7 & x8 & ~x5 & ~x6))) | (~x0 & x5 & x6 & ~x7 & ((x1 & ((x4 & x8) | (x3 & ~x4 & ~x8))) | (~x4 & x8 & ~x1 & ~x3)));
  assign z32 = (x4 & ((x2 & ((x1 & ((~x3 & ((~x0 & ((~x5 & ~x7 & x8) | (x7 & ~x8 & x5 & x6))) | (x7 & ((~x5 & x6 & x8) | (x0 & ~x6 & (~x5 | (x5 & x8))))) | (x5 & ~x7 & (~x6 | (x0 & x6 & x8))))) | (~x0 & ((x7 & ~x8 & ~x5 & ~x6) | (x3 & ((x7 & ~x8 & x5 & ~x6) | (~x5 & x6 & (~x7 ^ ~x8)))))))) | (~x1 & ((x3 & (x8 ? ((x5 & ~x6 & x7) | (x0 & (x5 ? ~x7 : (~x6 & x7)))) : (x0 ? ((~x5 & x6 & x7) | (~x6 & (~x7 | (x5 & x7)))) : (~x5 | (x5 & x6))))) | (~x3 & ((x5 & ((x6 & ~x7 & x8) | (x0 & (x8 ? x7 : x6)))) | (x7 & ~x8 & ~x0 & ~x6))) | (x6 & x7 & x8 & ~x0 & ~x5))) | (~x5 & x6 & ~x7 & x0 & ~x3))) | (~x2 & ((x1 & ((x5 & ((x7 & (x0 ? (~x6 & ~x8) : (x3 ? (x6 & x8) : ~x6))) | (x0 & ~x7 & (x3 ? (x6 & ~x8) : x8)))) | (x0 & ((~x3 & ((x6 & ~x7 & ~x8) | (~x5 & ~x6 & x8))) | (~x5 & x6 & x8 & (x7 | (x3 & ~x7))))))) | (~x1 & ((~x7 & (x0 ? (x3 ? (x5 & ~x8) : (~x5 & ~x6)) : (~x6 & (x3 ? ~x5 : (x5 & ~x8))))) | (~x3 & ((x7 & x8 & x5 & x6) | (~x5 & ((x7 & ~x8 & x0 & x6) | (~x0 & ~x6 & x8))))))) | (~x5 & ~x8 & ((x0 & x3 & ~x6 & x7) | (x6 & ~x7 & ~x0 & ~x3))))) | (~x5 & x7 & x8 & x0 & ~x1 & ~x3))) | (~x4 & ((x2 & ((x0 & (x5 ? (x6 ? (x1 ? (x7 & (~x8 | (x3 & x8))) : (x3 & ~x8)) : ((x8 & (x1 ? (~x3 | (x3 & ~x7)) : x3)) | (~x1 & ~x3 & ~x7))) : ((x3 & (x1 ? (~x8 & (~x6 ^ x7)) : (~x6 | (x6 & ~x7)))) | (x7 & (x1 ? x8 : (x6 & ~x8)))))) | (~x0 & ((x1 & ((x5 & ((~x3 & x7 & x8) | (~x7 & ~x8 & x3 & ~x6))) | (~x3 & x6 & ~x8) | (x8 & (x3 ? ((x6 & x7) | (~x5 & ~x6 & ~x7)) : (~x5 & ~x6))))) | (~x1 & x3 & x5 & x6 & x7) | (~x6 & ((~x3 & x5 & ~x7) | (~x1 & x7 & (x5 ? x8 : ~x3)))))) | (x1 & x3 & x6 & ~x7 & (x5 ^ ~x8)))) | (~x2 & ((x5 & ((~x0 & ((x3 & ~x6) | (x7 & ~x8 & x1 & ~x3))) | (x0 & ((~x6 & (x1 ? (~x8 & (~x3 | (x3 & x7))) : (~x3 & x8))) | (~x3 & x6 & (x7 ? x8 : ~x1)))) | (x1 & x3 & x6 & ~x7 & ~x8))) | (x7 & ((x3 & ((~x0 & (x1 ? (~x5 & ~x8) : x6)) | (~x6 & x8 & x0 & ~x1))) | (x1 & ((x0 & ((x6 & ~x8) | (~x3 & ~x6 & x8))) | (x6 & x8 & ~x0 & ~x5))))) | (~x5 & ((~x7 & ((x0 & ~x1 & (x3 ^ x8)) | (~x6 & ~x8 & x1 & ~x3))) | (~x0 & x1 & x3 & ~x6 & x8))) | (x6 & ~x7 & x8 & x0 & x1 & ~x3))) | (~x0 & ~x1 & ~x3 & ~x7 & x8 & x5 & x6))) | (x3 & ((~x6 & (x0 ? (x1 & ~x2 & (~x7 | (~x5 & x7 & x8))) : (~x1 & x2 & (x5 ? ~x8 : (x7 & x8))))) | (x0 & x5 & x6 & x8 & (x1 ? (~x2 & ~x7) : (x2 & x7))))) | (~x3 & ((x0 & ~x6 & ~x8 & ((~x1 & x5 & x7) | (x1 & x2 & ~x5 & ~x7))) | (~x7 & x8 & ~x5 & x6 & ~x0 & ~x1 & x2)));
  assign z33 = (x2 & ((x3 & ((x5 & (x8 ? (x6 ? (x0 ? (~x4 & x7) : (x1 ? (~x4 | (x4 & ~x7)) : (x4 & x7))) : (x0 ? (x1 ? (~x4 & ~x7) : (~x4 | (x4 & ~x7))) : (x4 & ~x7))) : ((x0 & ~x1 & ~x4 & x6) | (~x0 & x1 & x4 & ~x6 & x7)))) | (~x5 & ((x0 & ((~x4 & (x1 ? (x7 ? x6 : ~x8) : (~x6 | (x6 & ~x7)))) | (~x1 & x4 & ((~x6 & ~x7) | (x7 & x8) | (x6 & ~x8))))) | (x8 & ((x1 & ~x6 & ((~x4 & x7) | (~x0 & x4 & ~x7))) | (~x0 & x6 & (~x4 ^ ~x7)))) | (~x0 & x7 & ~x8 & (x1 ? (x4 & x6) : ~x4)))) | (~x0 & ~x4 & ~x7 & ~x8 & (~x1 ^ ~x6)))) | (x8 & ((~x0 & ((~x4 & ((x1 & ~x3 & ~x5 & x6) | (~x6 & ~x7 & ~x1 & x5))) | (~x3 & (x1 ? (~x7 & (x5 ? x6 : x4)) : (~x6 & x7 & (~x5 | (x4 & x5))))) | (~x1 & x4 & x5 & x6 & ~x7))) | (~x3 & ((x0 & ((~x4 & (x1 ? (x5 ? ~x6 : x7) : (~x5 & ~x7))) | (x4 & (x1 ? (x5 & (~x6 ^ ~x7)) : (x6 & x7))) | (x6 & ~x7 & ~x1 & x5))) | (x5 & ~x6 & ~x7 & x1 & x4))))) | (~x8 & ((~x3 & ((x5 & ((x0 & (x1 ? (x4 ? (~x6 & ~x7) : (x6 & x7)) : (x4 & x6))) | (~x6 & ((~x0 & x4 & ~x7) | (~x1 & ~x4 & x7))))) | (~x0 & ~x5 & ((~x1 & x6 & ~x7) | (x4 & ~x6 & x7))))) | (x6 & x7 & ((x4 & x5 & ~x0 & x1) | (x0 & ~x1 & ~x4 & ~x5))))) | (x0 & ~x3 & ((~x5 & ((x1 & ((~x6 & ~x7) | (x4 & x6 & x7))) | (x4 & (~x6 ^ ~x7)))) | (x5 & ~x6 & ~x7 & ~x1 & ~x4))))) | (~x2 & ((~x0 & ((((x6 & x7 & x3 & ~x4) | (~x6 & ~x7 & ~x3 & x4)) & (x1 ? (~x5 & ~x8) : (x5 & x8))) | (x8 & ((x1 & ~x3 & x4 & ~x5 & x6) | (~x6 & x7 & ~x4 & x5))) | (~x4 & ((~x6 & ((~x7 & (x1 ? (x5 ? ~x8 : x3) : x3)) | (~x1 & ~x3 & x5 & ~x8))) | (~x1 & x3 & x7 & (x5 ? ~x8 : x6)))) | (~x3 & x4 & ((~x8 & (x5 ? (x1 ? x7 : (x6 & ~x7)) : (x6 & x7))) | (~x1 & ~x5 & (~x6 | (x6 & ~x7))))))) | (x4 & ((x0 & ((x6 & (x1 ? (x7 ? (x5 ? (~x3 ^ x8) : x8) : ~x5) : ((~x3 & ~x5 & x7) | (~x7 & ~x8 & x3 & x5)))) | (~x6 & ((~x3 & ~x5 & x8) | (x5 & ((x3 & ~x7) | (x1 & (x3 ? (x7 & ~x8) : ~x7)))))) | (x1 & x3 & ~x5 & x7 & ~x8))) | (x5 & x6 & x8 & (~x1 ^ ~x7)))) | (x0 & (x1 ? ((~x6 & x8 & x3 & ~x5) | (~x3 & ((x7 & ((x5 & ((~x6 & ~x8) | (~x4 & x6 & x8))) | (~x4 & (x6 ^ x8)))) | (~x7 & x8 & ~x4 & x6)))) : (~x4 & ((~x7 & ~x8 & ~x5 & ~x6) | (x3 & (x6 ? (~x7 & ~x8) : (x7 & x8))))))) | (x1 & x3 & ~x4 & x5 & ~x6 & (~x7 ^ ~x8)))) | (x5 & ((~x4 & x6 & ((x1 & x3 & (x0 ? (~x7 ^ ~x8) : (~x7 & ~x8))) | (~x0 & ~x1 & ~x3 & ~x7 & x8))) | (x7 & ~x8 & x4 & ~x6 & x0 & ~x1 & ~x3))) | (~x1 & x3 & x4 & ~x5 & ~x6 & (x0 ? (x7 & ~x8) : (~x7 & x8)));
  assign z34 = (x2 & ((x1 & ((~x3 & (x5 ? ((~x8 & ((x6 & x7 & ~x0 & ~x4) | (~x6 & ~x7 & x0 & x4))) | (~x0 & ~x4 & (x7 ? x8 : x6)) | (x0 & x8 & ((~x6 & ~x7) | (x4 & (~x6 ^ ~x7))))) : ((x4 & ((~x6 & ~x7 & x8) | (x0 & (x7 | (x6 & ~x7))))) | (~x0 & ~x4 & (x6 | (~x6 & x8)))))) | (x3 & ((~x5 & ((~x0 & ((~x7 & x8 & ~x4 & ~x6) | (x4 & (x6 ? (~x7 & x8) : (x7 & ~x8))))) | (~x4 & ((x6 & (~x7 ^ x8)) | (x7 & x8 & x0 & ~x6))))) | (x0 & ~x4 & ((x6 & x7 & ~x8) | (x5 & x8 & (~x6 ^ x7)))) | (x6 & x7 & ~x8 & ~x0 & x4 & x5))) | (~x6 & ~x7 & ~x8 & x0 & ~x4 & ~x5))) | (~x1 & ((~x5 & (x0 ? ((x8 & (x3 ? ((~x6 & x7) | (x4 & (~x6 ^ x7))) : (~x4 & (~x6 | (x6 & ~x7))))) | (x6 & ~x7 & ~x8 & x3 & x4)) : (x3 ? (x4 & (~x6 ^ ~x7)) : (x6 ? (~x7 & x8) : x7)))) | (~x0 & ((x5 & ((x3 & ((x4 & (x6 ? x8 : ~x7)) | (~x7 & ~x8 & ~x4 & x6))) | (~x6 & x7 & (x8 | (x4 & ~x8))))) | (x6 & x7 & ~x8 & x3 & x4))) | (x0 & x4 & x7 & (x3 ? (~x6 & (~x8 | (x5 & x8))) : x8)))) | (~x0 & ~x3 & ((~x6 & ~x7 & ~x4 & x5) | (x6 & x7 & x8 & x4 & ~x5))))) | (~x1 & ((x3 & ((x4 & ((~x6 & (x0 ? ((x5 & ~x7 & x8) | (~x2 & ~x5 & x7)) : (~x5 & ~x7))) | (~x0 & x6 & (x5 ? (~x7 & ~x8) : (x7 & x8))))) | (~x0 & ~x4 & ((~x5 & ((x7 & x8) | (~x2 & ~x7 & (~x8 | (x6 & x8))))) | (x5 & ~x6 & ~x7) | (x7 & ((x6 & ~x8) | (x5 & (x6 ^ ~x8)))))))) | (~x3 & ((~x2 & (x0 ? ((~x5 & (x4 ? (~x8 & (~x6 ^ x7)) : (~x6 & ~x7))) | (x8 & ((x5 & x6 & x7) | (~x4 & (x6 ? ~x7 : x5))))) : ((~x5 & (x6 ? ~x7 : x4)) | (~x6 & ~x8 & ~x4 & x5)))) | (x5 & ((~x0 & ~x7 & (x4 ? ~x6 : (x6 & x8))) | (x0 & ~x4 & ~x6 & x7 & ~x8))))) | (~x7 & ~x8 & x5 & x6 & x0 & ~x2 & ~x4))) | (~x2 & ((x3 & ((x8 & ((~x0 & x1 & x4 & x5 & x6) | (x0 & ~x4 & ~x5 & ~x6 & ~x7))) | (x1 & ((~x7 & ((x0 & (x4 ? (~x5 | (x5 & x6 & ~x8)) : (~x6 & ~x8))) | (~x4 & x5 & (x6 ? ~x8 : ~x0)))) | (~x4 & ((x7 & ~x8 & x5 & ~x6) | (~x0 & ~x5 & (~x6 | (x6 & x7))))) | (x6 & x7 & ~x8 & x0 & ~x5))))) | (x1 & ((~x3 & (x0 ? ((~x6 & x7 & ~x8 & ~x4 & x5) | (x6 & ((x7 & x8 & ~x4 & x5) | (x4 & ~x8 & (~x7 | (x5 & x7)))))) : ((x4 & ((~x5 & x6 & x8) | (x7 & ~x8 & x5 & ~x6))) | (~x7 & ~x8 & ~x5 & ~x6)))) | (x0 & x4 & x5 & ~x7 & (~x6 | (x6 & x8))))) | (~x0 & x7 & ((~x6 & x8 & ~x4 & x5) | (~x3 & x4 & ~x5 & x6 & ~x8))) | (~x7 & x8 & ~x5 & x6 & x0 & ~x3 & x4))) | (x3 & ~x4 & x0 & x1 & ~x7 & x8 & x5 & x6);
  assign z35 = (x7 & ((x2 & ((x5 & (x0 ? (x3 ? ((~x4 & x6 & ~x8) | (~x6 & x8 & ~x1 & x4)) : (x1 ? (~x4 & (x6 ^ x8)) : (~x8 & (~x6 | (x4 & x6))))) : ((~x1 & x3 & (x4 ? (~x6 | (x6 & ~x8)) : (~x8 | (x6 & x8)))) | (~x6 & x8 & ~x3 & ~x4)))) | (~x5 & ((~x1 & ((~x4 & (x0 ? (x3 ? ~x8 : (~x6 & x8)) : ~x6)) | (~x0 & x4 & (x3 ^ x8)))) | (~x0 & x1 & x3 & (x4 ? (~x6 & ~x8) : (x6 & x8))))) | (x4 & ~x6 & ~x8 & x0 & ~x1 & x3))) | (x4 & ((~x2 & (x0 ? (x1 ? ((x5 & ~x6 & ~x8) | (x6 & x8 & x3 & ~x5)) : (~x5 & (x3 ? ~x6 : (x6 & ~x8)))) : ((x1 & x5 & (x3 ? (x6 & x8) : ~x6)) | (x6 & x8 & ~x1 & ~x3)))) | (~x0 & ~x1 & x8 & (x3 ? (~x5 & x6) : (x5 & ~x6))))) | (~x2 & (x0 ? ((~x3 & ((~x6 & x8 & x1 & ~x4) | (~x1 & x5 & (x8 ? x6 : ~x4)))) | (x1 & ((~x4 & x6 & ~x8) | (~x6 & x8 & x3 & ~x5)))) : (x1 & ~x4 & (x3 ? (~x5 & ~x8) : (x5 ? ~x8 : (x6 & x8)))))))) | (x2 & ((x8 & (x1 ? ((~x4 & (x0 ? ((x3 & x5 & x6) | (~x6 & ~x7 & ~x3 & ~x5)) : (~x5 & ~x6 & (~x3 | (x3 & ~x7))))) | (~x0 & x4 & ~x5 & ~x7 & (~x3 | (x3 & x6)))) : ((~x7 & (x0 ? ((~x4 & x5 & ~x6) | (~x3 & x4 & x6)) : (x3 ? (x6 ? x4 : x5) : (x5 ? x4 : x6)))) | (~x0 & x3 & x4 & ~x5 & ~x6)))) | (~x7 & ((~x1 & ((~x3 & x4 & ~x5 & x6 & ~x8) | (x3 & ((x6 & ~x8 & ~x4 & x5) | (x0 & ~x6 & (x4 ? (x5 & ~x8) : ~x5)))))) | (~x0 & ~x4 & ((~x3 & x5 & ~x6) | (x1 & x6 & ~x8 & (~x3 ^ ~x5)))))) | (~x0 & x1 & ~x3 & x6 & ~x8 & ~x4 & ~x5))) | (~x2 & ((~x0 & (x3 ? ((x1 & ~x4 & ~x5 & ~x6 & x8) | (x6 & ~x7 & ~x8 & ~x1 & x4 & x5)) : (~x7 & ((~x1 & x4 & x5 & ~x6 & ~x8) | (~x5 & ((~x6 & x8 & ~x1 & x4) | (x1 & ~x8 & (~x4 ^ x6)))))))) | (x0 & ((~x7 & ((~x3 & ((x8 & (x1 ? (x4 ? x5 : x6) : (~x4 & ~x5))) | (~x1 & ~x8 & (x4 ? (~x5 & ~x6) : x6)))) | (x1 & x3 & ~x4 & ((~x6 & ~x8) | (x5 & (x6 ^ x8)))))) | (~x6 & ((x1 & x4 & ~x5 & (x3 ^ x8)) | (~x1 & ~x3 & ~x4 & x5 & x8))))) | (~x7 & x8 & x5 & x6 & ~x1 & ~x3 & ~x4)));
  assign z36 = (x1 & ((~x2 & ((x3 & ((x5 & ((x7 & ((~x8 & (x0 ? (~x4 ^ ~x6) : (~x4 & ~x6))) | (x6 & x8 & ~x0 & x4))) | (~x4 & ~x7 & (x0 ? (~x6 & x8) : (x6 & ~x8))))) | (~x5 & ((x0 & ((~x6 & ~x7 & ~x8) | (x7 & ((~x6 & x8) | (x4 & (~x8 | (x6 & x8))))))) | (~x4 & ((x6 & x7 & ~x8) | (~x0 & ~x6 & ~x7))))) | (x6 & ~x7 & ~x8 & x0 & x4))) | (~x3 & ((x0 & ((x4 & ((x7 & ~x8 & x5 & x6) | (~x5 & ~x6 & x8))) | (~x4 & x7 & (x6 ^ x8)) | (~x7 & ((x6 & x8) | (x5 & ~x6 & ~x8))))) | (x4 & ((x7 & ~x8 & x5 & ~x6) | (~x0 & ((x6 & x7 & ~x8) | (~x5 & (x8 ? x6 : ~x7)))))))) | (x6 & ~x7 & x8 & ~x0 & x4 & x5))) | (x2 & ((x7 & (x3 ? ((~x5 & ((x0 & ~x4 & (x8 | (x6 & ~x8))) | (~x6 & ~x8 & ~x0 & x4))) | (x5 & x6 & ~x8 & ~x0 & x4)) : ((x0 & (x4 ? (~x5 | (x5 & ~x6 & x8)) : (x5 & ~x6))) | (~x4 & x5 & (x8 ? ~x0 : x6))))) | (~x7 & (x3 ? (~x5 & ((~x0 & x8 & (~x4 ^ x6)) | (~x4 & ~x8 & (x6 | (x0 & ~x6))))) : (x4 ? ((~x5 & ~x6 & x8) | (x0 & (x5 ? (~x6 & ~x8) : x6))) : ((~x0 & x5) | (~x6 & x8 & x0 & ~x5))))) | (~x0 & ~x3 & ~x4 & ~x5 & (x6 | (~x6 & x8))))) | (x0 & ~x3 & x4 & ~x7 & x8 & x5 & ~x6))) | (~x1 & ((x0 & ((x4 & (x3 ? (x5 ? ((~x6 & (x2 ? (~x8 | (x7 & x8)) : (~x7 & x8))) | (x7 & ~x8 & ~x2 & x6)) : ((~x6 & x7 & ~x8) | (x2 & x8 & (~x6 ^ x7)))) : ((x2 & ((x5 & x6 & (~x7 ^ ~x8)) | (~x6 & x7 & ~x8))) | (~x5 & ~x8 & ((~x6 & ~x7) | (~x2 & x6 & x7)))))) | (~x3 & ((x5 & ((x7 & x8 & ~x2 & x6) | (~x4 & (x2 ? (x6 ? (x7 & x8) : ~x8) : ~x6)))) | (~x4 & ((x6 & ~x7 & x8) | (x2 & ~x5 & (x6 ? (x7 & ~x8) : x8)))))) | (~x4 & ((x3 & ~x5 & ~x6 & ~x7 & x8) | (~x8 & ((x6 & (x2 ? (x3 & (~x7 | (x5 & x7))) : (x5 & ~x7))) | (~x5 & ~x6 & x2 & x3))))))) | (~x0 & ((x4 & ((x2 & x8 & ((x5 & x6 & ~x7) | (x3 & (x5 ? (x6 & x7) : ~x7)))) | (~x7 & ((x5 & ((~x3 & ~x6) | (~x2 & x6 & ~x8))) | (~x6 & ~x8 & x3 & ~x5))) | (~x2 & ~x3 & ~x5 & (x6 | (~x6 & ~x8))))) | (x5 & ((~x8 & (x2 ? (x3 ? (x6 & ~x7) : (~x6 & x7)) : (~x4 & (x3 ? x7 : ~x6)))) | (x2 & x3 & ~x6 & (~x7 | (~x4 & x7 & x8))))) | (x3 & ((~x2 & ((x7 & x8 & ~x5 & x6) | (~x7 & ~x8 & ~x4 & ~x6))) | (x2 & ~x4 & ~x5 & x7 & ~x8))))) | (x2 & x4 & ((~x3 & ((~x5 & x6 & ~x7) | (x7 & x8 & x5 & ~x6))) | (x6 & ~x7 & ~x8 & x3 & ~x5))) | (~x2 & ~x3 & ~x4 & ~x5 & ~x6 & ~x7))) | (x8 & ((~x0 & ((x7 & ((x5 & ~x6 & ~x2 & ~x3) | (x2 & ~x5 & x6 & (x3 ^ x4)))) | (~x2 & x3 & ~x4 & x5 & ~x6))) | (~x6 & ~x7 & ~x4 & x5 & x0 & x2 & x3)));
  assign z37 = (~x1 & ((~x5 & ((~x2 & ((~x6 & ((x0 & (x3 ? ~x4 : (x4 & ~x7))) | (x4 & x7 & ~x0 & ~x3))) | (~x0 & ((~x4 & (x3 ? (x8 ? ~x7 : x6) : (x6 & ~x7))) | (x6 & ~x8 & ~x3 & x4))) | (x6 & x7 & x8 & ~x3 & x4))) | (x2 & (x7 ? ((x0 & x6 & ((x4 & x8) | (~x3 & ~x4 & ~x8))) | (~x0 & x4 & (x8 ? x3 : ~x6)) | (~x4 & ~x6 & (x3 ^ x8))) : ((x3 & x4 & ~x8) | (~x4 & (x0 ? (x3 ? (~x6 | (x6 & x8)) : x8) : (x6 & ~x8)))))) | (~x6 & ~x7 & x8 & ~x0 & x3 & x4))) | (x5 & ((x0 & ((x4 & ((~x6 & ~x7 & ~x2 & x3) | (x6 & ~x8 & x2 & ~x3))) | (~x4 & ((x7 & (x2 ? (x3 ? x6 : (~x6 & ~x8)) : (~x6 & (~x3 | (x3 & x8))))) | (x6 & ~x7 & (x2 ? (~x3 & x8) : ~x8)))) | (x6 & x7 & x8 & ~x2 & ~x3))) | (~x0 & (x7 ? ((~x2 & x8 & (x3 ? ~x4 : ~x6)) | (x6 & ~x8 & x3 & ~x4)) : ((x2 & (x3 ? ~x6 : (~x4 & x8))) | (x4 & (x3 ? (x6 & ~x8) : ~x6))))) | (x2 & ((~x6 & x7 & ((x4 & x8) | (x3 & (x4 ^ x8)))) | (x6 & ~x7 & ~x8 & x3 & ~x4))))) | (~x0 & x2 & x3 & x4 & x6 & (~x7 ^ ~x8)) | (x0 & ~x2 & ~x3 & ~x4 & ~x6 & ~x7))) | (x1 & (x0 ? ((x4 & (x2 ? (~x3 & (((~x7 | (x7 & x8)) & (~x5 ^ ~x6)) | (~x5 & ~x6 & x7) | (~x7 & x8 & x5 & x6))) : ((x6 & (x3 ? (x5 ? (~x7 & x8) : x7) : (~x7 & x8))) | (~x7 & x8 & x5 & ~x6) | (~x3 & (x5 ? (x7 & ~x8) : (~x6 & x8)))))) | (~x3 & (x2 ? (~x5 & ((~x4 & x7 & x8) | (~x6 & ~x7 & ~x8))) : (~x4 & (x6 ? (x7 & ~x8) : (~x7 ^ x8))))) | (~x2 & x3 & ~x4 & x5 & x7 & ~x8)) : (x4 ? (x6 & ((x2 & (x5 ? (x7 & ~x8) : (x3 ? (~x7 ^ ~x8) : x7))) | (~x2 & ~x3 & ~x5 & ~x7 & ~x8))) : ((~x2 & ((~x6 & (x3 ? (x5 ? (~x7 & ~x8) : x8) : (x5 & ~x8))) | (~x5 & x7 & (x8 ? x6 : x3)))) | (x2 & ((~x3 & x5 & ~x7) | (x8 & ((~x3 & x5 & x7) | (x6 & (x3 ? (x7 | (x5 & ~x7)) : ~x5)))))) | (x6 & x7 & ~x8 & ~x3 & x5))))) | (x0 & ~x2 & x6 & ~x7 & (x3 ? (x4 & (~x5 ^ ~x8)) : (~x4 & x8)));
  assign z38 = (x8 & ((x1 & (((x3 ^ x4) & ((x0 & ((~x6 & x7 & x2 & ~x5) | (x6 & ~x7 & ~x2 & x5))) | (~x0 & ~x2 & x5 & ~x6 & x7))) | (~x5 & (x3 ? ((x2 & ((~x4 & x6 & x7) | (~x0 & ~x7 & (~x4 ^ x6)))) | (~x6 & ~x7 & x0 & ~x2)) : ((x4 & ((x6 & (x0 ? (~x2 ^ ~x7) : x7)) | (~x0 & x2 & ~x7))) | (x0 & ~x4 & (x6 ? (x2 ^ ~x7) : x7))))) | (x5 & ((x0 & ((~x4 & ((x2 & ~x6 & (x3 ^ x7)) | (x6 & x7 & ~x2 & ~x3))) | (~x6 & ~x7 & ~x2 & ~x3))) | (~x0 & x2 & ~x3 & ~x4 & x7))))) | (~x1 & ((x6 & ((x5 & ((x2 & (x0 ? (x7 & (~x4 | (x3 & x4))) : (~x7 & (~x3 | (x3 & x4))))) | (x0 & ~x3 & ((~x2 & ~x4 & ~x7) | (x4 & x7))))) | (~x0 & ((~x2 & ~x5 & (x3 ? (x4 & x7) : ~x7)) | (x2 & x3 & ~x4 & x7))) | (x4 & ~x5 & ~x7 & x0 & ~x2 & ~x3))) | (~x6 & ((~x4 & ((x5 & (x0 ? (x2 ? x3 : x7) : (x3 & ~x7))) | (~x5 & x7 & ~x2 & x3))) | (x2 & x5 & (x0 ? (x4 & x7) : (x7 ? x3 : x4))))) | (x0 & ~x5 & ((x2 & ~x4 & ~x7) | (~x2 & ~x3 & x4 & x7))))) | (x0 & ~x2 & x3 & ~x6 & x7 & x4 & ~x5))) | (~x8 & ((~x1 & ((x3 & ((~x7 & (x0 ? ((~x2 & (x4 ? x5 : x6)) | (~x5 & ~x6 & x2 & x4)) : ((x4 & x5 & x6) | (x2 & (x6 ? ~x4 : x5))))) | (~x6 & ((x7 & ((x0 & x5 & (x2 ^ ~x4)) | (x2 & ~x4 & ~x5))) | (x0 & ~x2 & ~x4 & ~x5))))) | (~x3 & ((~x7 & (x0 ? ((x4 & ~x5 & ~x6) | (~x2 & ~x4 & x5)) : ((x4 & x5 & ~x6) | (~x2 & ~x4 & ~x5)))) | (x0 & x7 & ((x4 & ((x5 & ~x6) | (~x2 & ~x5 & x6))) | (~x5 & x6 & x2 & ~x4))))) | (~x0 & ~x4 & x5 & ~x6 & x7))) | (x1 & ((x7 & ((x2 & ((~x3 & x6 & (x0 ? (~x4 ^ ~x5) : ~x4)) | (~x0 & x3 & x4 & ~x5))) | (x0 & ~x2 & ((~x5 & x6 & x3 & ~x4) | (~x3 & (x6 ? ~x4 : x5)))))) | (~x2 & ((~x7 & ((~x4 & (x0 ? (~x5 & ~x6) : (x5 & (~x6 | (x3 & x6))))) | (x0 & x3 & x4 & (x6 | (x5 & ~x6))))) | (~x0 & x3 & ~x4 & ~x5 & ~x6))) | (~x4 & ~x5 & ~x7 & x0 & x2 & x3))) | (~x5 & x7 & ((~x0 & ~x2 & x3 & ~x4 & x6) | (x0 & x2 & ~x3 & x4 & ~x6))))) | (x2 & ((~x7 & ((~x3 & ((x4 & ((x0 & (x1 ? (~x5 & ~x6) : (x5 & x6))) | (x1 & x5 & ~x6))) | (~x0 & x1 & ~x4 & x6))) | (~x0 & ~x1 & x3 & x4 & ~x5))) | (x0 & ~x1 & x3 & x6 & x7 & x4 & ~x5))) | (~x0 & ~x1 & ~x3 & ~x6 & x7 & x4 & ~x5);
  assign z39 = (x4 & ((x2 & (x1 ? ((~x0 & ((~x7 & x8 & x5 & x6) | (x3 & ((x7 & ~x8 & x5 & x6) | (~x6 & ~x7 & x8))))) | (~x3 & ((~x7 & ((x5 & ~x6 & ~x8) | (x0 & (x5 ? (x6 & x8) : ~x6)))) | (~x5 & ((x6 & x7 & x8) | (x0 & (x6 ? ~x8 : (x7 & x8)))))))) : (x5 ? ((x0 & (x3 ? (x6 ? (x7 & ~x8) : (~x7 ^ x8)) : ((x7 & x8) | (x6 & ~x7 & ~x8)))) | (x3 & ((x6 & x7 & x8) | (~x0 & (~x7 ^ ~x8)))) | (~x7 & ~x8 & ~x0 & ~x6)) : ((x3 & (x0 ? (x7 ? x6 : ~x8) : (x6 | (~x6 & ~x8)))) | (x6 & ~x7 & x8 & x0 & ~x3))))) | (~x1 & (x0 ? (~x2 & ((x3 & (x5 ? (x6 ? (x7 & x8) : ~x7) : (~x6 & x7))) | (~x3 & ~x5 & ~x6 & ~x7 & ~x8))) : ((~x7 & ((x5 & ~x6 & ~x2 & ~x3) | (x3 & (x5 ? (x6 & ~x8) : (~x6 & x8))))) | (~x2 & ~x3 & (x5 ? (x7 & x8) : (x6 ? x8 : (x7 & ~x8))))))) | (~x2 & ((x1 & ((~x3 & (x0 ? ((~x7 & x8 & ~x5 & x6) | (x5 & ~x8)) : (x5 ? (~x6 & x7) : (~x7 & ~x8)))) | (x0 & x3 & (x5 ? (~x6 & x7) : (~x7 & (~x6 | (x6 & ~x8))))))) | (x0 & x6 & ((~x7 & ~x8 & x3 & x5) | (x7 & x8 & ~x3 & ~x5))))) | (x7 & ~x8 & ~x5 & x6 & ~x0 & x1 & ~x3))) | (~x4 & ((x0 & ((~x7 & ((x3 & ((~x5 & ((~x1 & ((~x6 & ~x8) | (x2 & x6 & x8))) | (~x6 & ~x8 & x1 & x2))) | (x1 & ((~x2 & ~x6) | (x5 & ((x6 & ~x8) | (x2 & ~x6 & x8))))))) | (~x2 & ~x3 & (x1 ? (x6 & x8) : (~x6 | (x6 & ~x8)))))) | (x7 & (x1 ? ((x6 & (x2 ? (x5 ? (~x8 | (x3 & x8)) : x8) : (x3 ? (~x5 & ~x8) : (x5 & x8)))) | (x2 & x3 & ~x5 & ~x6 & x8)) : ((x8 & (x2 ? (x3 ? x5 : (~x5 & ~x6)) : (x3 & ~x6))) | (~x2 & ~x3 & x5 & x6)))) | (x1 & ~x2 & ~x3 & ~x6 & (x5 | (~x5 & x8))))) | (x5 & ((~x0 & (x1 ? ((~x8 & (x2 ? (~x7 & (x6 | (x3 & ~x6))) : (x3 ? ~x6 : x7))) | (x2 & ~x3 & x8 & (~x6 ^ x7))) : ((x7 & ((x3 & x6 & x8) | (~x2 & ~x6 & ~x8))) | (x3 & ~x6 & (x8 ? x2 : ~x7))))) | (x2 & x3 & x6 & (x1 ? (~x7 & x8) : ~x8)))) | (~x0 & ((x1 & ((x2 & ((x7 & ~x8 & ~x3 & x6) | (~x6 & ~x7 & x3 & ~x5))) | (~x3 & ((x7 & x8 & ~x5 & x6) | (~x7 & ~x8 & ~x2 & ~x6))))) | (x3 & ~x5 & x7 & ((~x6 & x8) | (~x2 & x6 & ~x8))))) | (x1 & x2 & ~x5 & ((x7 & x8 & ~x3 & ~x6) | (~x7 & ~x8 & x3 & x6))))) | (~x8 & ((x0 & ~x1 & x2 & ~x5 & x7 & (~x3 ^ ~x6)) | (~x0 & x1 & ~x2 & x6 & ~x7 & x3 & x5))) | (x2 & ~x3 & x8 & ((x5 & ((x0 & (x1 ? (~x6 & x7) : (x6 & ~x7))) | (~x6 & ~x7 & ~x0 & ~x1))) | (~x0 & ~x5 & (x1 ? (x6 & ~x7) : (~x6 & x7)))));
endmodule