module pla__b12 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14,
    z0, z1, z2, z3, z4, z5, z6, z7, z8  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14;
  output z0, z1, z2, z3, z4, z5, z6, z7, z8;
  assign z0 = ~x00 & ((x01 & (((~x04 | x05) & (x02 | x03)) | (~x02 & x03))) | (x02 & x03 & ~x04));
  assign z1 = ~x00 & ((x02 & (x03 | x04) & (~x01 | ~x05 | ~x06)) | (x01 & x03 & (~x02 | ~x05 | ~x06)));
  assign z2 = ((~x00 | (~x07 & ~x08)) & (x02 | (~x01 & ~x03 & (x09 | x10)))) | (~x01 & ((~x00 & (x07 ? ~x03 : (x09 & ~x10))) | (~x07 & ~x08 & x09 & ~x10)));
  assign z3 = (~x07 | ~x11) & (x00 | ~x12);
  assign z4 = ((~x07 | ~x11) & (~x00 | ~x08 | ~x09)) | (x07 & ~x11);
  assign z5 = x12 | ~x13 | x10 | x00 | x07;
  assign z6 = ~x07 & ~x10 & (((x01 | x02 | (~x03 & x09) | (x03 & ~x09)) & ((~x08 & (x00 | ~x14)) | (~x00 & ~x14))) | ((~x00 | ~x08) & (((x03 ^ x09) & (~x01 | ~x02)) | (~x01 & x02) | (x01 & ~x02))));
  assign z7 = (x09 & (~x08 | (~x01 & ~x02 & x03))) | (~x08 & (x01 | x02 | ~x03)) | x07 | x10;
  assign z8 = ((~x00 | x09) & (x01 | x02 | ~x03 | x12)) | x07 | x10 | (~x00 & ~x09);
endmodule