module pla__x7dn ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55,
    x56, x57, x58, x59, x60, x61, x62, x63, x64, x65,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54,
    x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14;
  assign z00 = (x00 | x01) & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x02 : x05)) | (x05 & ~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))));
  assign z01 = ((x04 | (x06 & x08 & x09 & ~x10)) & (((x00 | x01) & (x03 ? x11 : x12)) | (~x00 & ~x01 & ((x13 & (~x14 | (~x03 & x14 & ~x15))) | (x03 & x16))))) | (~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09)) & ((x12 & (x00 | x01)) | (~x00 & ~x01 & x13)));
  assign z02 = ((x04 | (x06 & x08 & x09 & ~x10)) & (((x00 | x01) & (x03 ? x17 : x18)) | (~x00 & ~x01 & ((x19 & (~x14 | (~x03 & x14 & ~x15))) | (x03 & x20))))) | (~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09)) & ((x18 & (x00 | x01)) | (~x00 & ~x01 & x19)));
  assign z03 = ((x04 | (x06 & x08 & x09 & ~x10)) & (((x00 | x01) & (x03 ? x21 : x22)) | (~x00 & ~x01 & ((x23 & (~x14 | (~x03 & x14 & ~x15))) | (x03 & x24))))) | (~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09)) & ((x22 & (x00 | x01)) | (~x00 & ~x01 & x23)));
  assign z04 = ((x04 | (x06 & x08 & x09 & ~x10)) & (((x00 | x01) & (x03 ? x25 : x26)) | (~x00 & ~x01 & ((x27 & (~x14 | (~x03 & x14 & ~x15))) | (x03 & x28))))) | (~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09)) & ((x26 & (x00 | x01)) | (~x00 & ~x01 & x27)));
  assign z05 = ((x04 | (x06 & x08 & x09 & ~x10)) & (((x00 | x01) & (x03 ? x29 : x30)) | (~x00 & ~x01 & ((x31 & (~x14 | (~x03 & x14 & ~x15))) | (x03 & x32))))) | (~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09)) & ((x30 & (x00 | x01)) | (~x00 & ~x01 & x31)));
  assign z06 = ((x04 | (x06 & x08 & x09 & ~x10)) & (((x00 | x01) & (x03 ? x33 : x34)) | (~x00 & ~x01 & ((x35 & (~x14 | (~x03 & x14 & ~x15))) | (x03 & x36))))) | (~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09)) & ((x34 & (x00 | x01)) | (~x00 & ~x01 & x35)));
  assign z07 = ((x04 | (x06 & x08 & x09 & ~x10)) & (((x00 | x01) & (x03 ? x37 : x38)) | (~x00 & ~x01 & (x03 ? x02 : x05)))) | (~x06 & (x07 ? (x09 & ~x10) : (~x08 ^ x09)) & ((x38 & (x00 | x01)) | (~x00 & ~x01 & x05)));
  assign z08 = (~x00 & ~x01 & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x11 : x12)) | (~x06 & x12 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))))) | ((x00 | x01) & ((~x06 & ((x09 & (x07 ? (~x10 & (x39 ? (x52 ? (~x45 | ~x46 | ~x47 | ~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x45 | x46 | x47 | x48 | x49 | x50 | x51)))) : ((x45 & x46 & x47 & x48 & x49 & x50 & x51 & x52) | (~x45 & ~x46 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & x53)))) : (x08 & x44))) | (~x07 & ~x08 & ~x09 & ((x41 & ~x43 & (x42 ? x39 : x44)) | (x40 & ~x42 & x43))))) | (x06 & x08 & x09 & ~x10 & (x07 ? x39 : (x39 ? (x52 ? (~x45 | ~x46 | ~x47 | ~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x45 | x46 | x47 | x48 | x49 | x50 | x51)))) : ((x45 & x46 & x47 & x48 & x49 & x50 & x51 & x52) | (~x45 & ~x46 & ~x47 & ~x48 & ~x49 & ~x50 & ~x51 & ~x52 & x53))))) | (x04 & x39)));
  assign z09 = (~x00 & ~x01 & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x17 : x18)) | (~x06 & x18 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))))) | ((x00 | x01) & ((~x06 & ((x09 & (x07 ? (~x10 & (x45 ? (x52 ? (~x46 | ~x47 | ~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x46 | x47 | x48 | x49 | x50 | x51)))) : ((x49 & x50 & x51 & x52 & x46 & x47 & x48) | (~x46 & ~x47 & ~x48 & ~x49 & ~x52 & x53 & ~x50 & ~x51)))) : (x08 & (x55 | (x03 & x10 & x56))))) | (~x07 & ~x08 & ~x09 & ((x41 & ~x43 & (x42 ? x45 : x55)) | (~x42 & x43 & x54))))) | (x06 & x08 & x09 & ~x10 & (x07 ? x45 : (x45 ? (x52 ? (~x46 | ~x47 | ~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x46 | x47 | x48 | x49 | x50 | x51)))) : ((x49 & x50 & x51 & x52 & x46 & x47 & x48) | (~x46 & ~x47 & ~x48 & ~x49 & ~x52 & x53 & ~x50 & ~x51))))) | (x04 & x45)));
  assign z10 = (~x00 & ~x01 & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x21 : x22)) | (~x06 & x22 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))))) | ((x00 | x01) & ((~x06 & (x07 ? (x09 & ~x10 & (x46 ? (x52 ? (~x47 | ~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x47 | x48 | x49 | x50 | x51)))) : ((x47 & x48 & x49 & x50 & x51 & x52) | (~x52 & x53 & ~x50 & ~x51 & ~x47 & ~x48 & ~x49)))) : ((x16 & ((x08 & x09) | (~x08 & ~x09 & x41 & ~x42 & ~x43))) | (~x08 & ~x09 & ((x13 & ~x42 & x43) | (x41 & x42 & ~x43 & x46)))))) | (x06 & x08 & x09 & ~x10 & (x07 ? x46 : (x46 ? (x52 ? (~x47 | ~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x47 | x48 | x49 | x50 | x51)))) : ((x47 & x48 & x49 & x50 & x51 & x52) | (~x52 & x53 & ~x50 & ~x51 & ~x47 & ~x48 & ~x49))))) | (x04 & x46)));
  assign z11 = (~x00 & ~x01 & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x25 : x26)) | (~x06 & x26 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))))) | ((x00 | x01) & ((~x06 & (x07 ? (x09 & ~x10 & (x47 ? (x52 ? (~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x48 | x49 | x50 | x51)))) : ((x48 & x49 & x50 & x51 & x52) | (~x51 & ~x52 & x53 & ~x48 & ~x49 & ~x50)))) : ((x20 & ((x08 & x09) | (~x08 & ~x09 & x41 & ~x42 & ~x43))) | (~x08 & ~x09 & ((x19 & ~x42 & x43) | (x41 & x42 & ~x43 & x47)))))) | (x06 & x08 & x09 & ~x10 & (x07 ? x47 : (x47 ? (x52 ? (~x48 | ~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x48 | x49 | x50 | x51)))) : ((x48 & x49 & x50 & x51 & x52) | (~x51 & ~x52 & x53 & ~x48 & ~x49 & ~x50))))) | (x04 & x47)));
  assign z12 = (~x00 & ~x01 & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x29 : x30)) | (~x06 & x30 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))))) | ((x00 | x01) & ((~x06 & (x07 ? (x09 & ~x10 & (x48 ? (x52 ? (~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x49 | x50 | x51)))) : ((x49 & x50 & x51 & x52) | (~x49 & ~x50 & ~x51 & ~x52 & x53)))) : ((x24 & ((x08 & x09) | (~x08 & ~x09 & x41 & ~x42 & ~x43))) | (~x08 & ~x09 & ((x23 & ~x42 & x43) | (x41 & x42 & ~x43 & x48)))))) | (x06 & x08 & x09 & ~x10 & (x07 ? x48 : (x48 ? (x52 ? (~x49 | ~x50 | ~x51) : (~x53 | (x53 & (x49 | x50 | x51)))) : ((x49 & x50 & x51 & x52) | (~x49 & ~x50 & ~x51 & ~x52 & x53))))) | (x04 & x48)));
  assign z13 = (~x00 & ~x01 & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x33 : x34)) | (~x06 & x34 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))))) | ((x00 | x01) & ((~x06 & (x07 ? (x09 & ~x10 & (x49 ? (x52 ? (~x50 | ~x51) : (~x53 | (x53 & (x50 | x51)))) : ((~x52 & x53 & ~x50 & ~x51) | (x50 & x51 & x52)))) : ((x28 & ((x08 & x09) | (~x08 & ~x09 & x41 & ~x42 & ~x43))) | (~x08 & ~x09 & ((x41 & x42 & ((~x43 & x49) | (x43 & x57 & x58 & ~x59 & ~x60 & ~x61 & ~x62 & ~x63))) | (x27 & ~x42 & x43)))))) | (x06 & x08 & x09 & ~x10 & (x07 ? x49 : (x49 ? (x52 ? (~x50 | ~x51) : (~x53 | (x53 & (x50 | x51)))) : ((~x52 & x53 & ~x50 & ~x51) | (x50 & x51 & x52))))) | (x04 & x49)));
  assign z14 = (~x00 & ~x01 & (((x04 | (x06 & x08 & x09 & ~x10)) & (x03 ? x37 : x38)) | (~x06 & x38 & (x07 ? (x09 & ~x10) : (~x08 ^ x09))))) | ((x00 | x01) & ((~x06 & (x07 ? (x09 & ~x10 & (x50 ? (x52 ? ~x51 : (~x53 | (x51 & x53))) : (x51 ? x52 : (~x52 & x53)))) : ((x32 & ((x08 & x09) | (~x08 & ~x09 & x41 & ~x42 & ~x43))) | (~x08 & ~x09 & ((x41 & x42 & (x43 ? (~x59 & ~x60 & ~x61 & ~x62 & (x58 ? (~x63 & x65) : (x63 & x64))) : x50)) | (x31 & ~x42 & x43)))))) | (x06 & x08 & x09 & ~x10 & (x07 ? x50 : (x50 ? (x52 ? ~x51 : (~x53 | (x51 & x53))) : (x51 ? x52 : (~x52 & x53))))) | (x04 & x50)));
endmodule