module pla__x6dn ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38,
    z0, z1, z2, z3, z4  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38;
  output z0, z1, z2, z3, z4;
  assign z0 = x01 & ((~x05 & ((~x00 & (x03 ? (x04 & (x02 ? ~x14 : (x14 & x19 & x26 & (~x22 | ~x23) & (~x27 | ~x28)))) : (x04 ? (~x14 & (x02 ? (x17 ? ~x13 : ((~x22 | ~x23) & (~x21 | (x18 & x19 & ~x20)))) : x16)) : (x02 ? (x14 & ((x16 & (~x17 | ~x19)) | (~x16 & (x17 | x19)) | (~x17 & x19) | ~x25 | (x17 & ~x19))) : (x06 & (~x07 | (x07 & ((~x08 & (x09 | (~x09 & ~x10 & ~x11 & x12))) | (x10 & ~x11 & ~x13 & (x08 | ~x09)))))))))) | (~x14 & ((x00 & (x02 ? (~x03 | (x03 & (x22 | x23 | (~x22 & ~x23)))) : (x03 ^ x04))) | (~x02 & x03 & x04 & (~x21 | (x17 & ~x20))))) | (x00 & ~x02 & x03 & x14))) | (x02 & (x03 ? (((x22 | x23) & ((x00 & (x04 ? (x05 & ~x14) : x14)) | (~x00 & x04 & x05 & ~x13 & ~x14 & x17))) | (x00 & ((x04 & x05 & (x14 | (~x14 & ~x22 & ~x23))) | (~x22 & ~x23 & ~x04 & x14))) | (~x04 & x05 & ~x14 & ~x17 & x18 & ~x20)) : ((x00 & ~x04 & x14) | (~x00 & x04 & x05 & ~x14 & x23 & ~x24)))) | (x00 & ((~x14 & (x03 ? (x04 ? ~x02 : x05) : (x04 & x05))) | (~x02 & ~x03 & (~x04 | (x04 & x14))))));
  assign z1 = x01 & ((~x05 & ((~x00 & (x02 ? (~x03 & (x04 ? (~x14 & ~x17 & (~x22 | ~x23) & (~x21 | (x18 & x19 & ~x20))) : (x14 & ((x16 & (~x17 | ~x19)) | (~x16 & (x17 | x19)) | (~x17 & x19) | ~x25 | (x17 & ~x19))))) : (x03 ? ((x04 & (x14 ? ((~x27 | ~x28) & ((x22 & x23) | (x19 & x26 & (~x22 | ~x23)))) : (x21 & (~x17 | x20) & (~x34 | (x19 & x34))))) | (x27 & x28 & x14 & x19)) : (x04 ? (~x14 & x16) : (x06 & (~x07 | (x07 & ((x10 & ((x08 & (x11 | (~x09 & ~x11 & x13))) | (~x09 & x11))) | (x09 & (~x08 | (x08 & (~x10 | (~x11 & x13))))))))))))) | (x00 & ~x02 & x03 & x14) | (~x14 & ((~x02 & ((x00 & (x03 ^ x04)) | (x03 & x04 & (~x21 | (x17 & ~x20))) | (~x03 & ~x04 & x29 & x30 & x31 & ~x32 & x33))) | (x00 & x02 & (~x03 | (x03 & (x22 | x23 | (~x22 & ~x23))))))))) | (x00 & (x03 ? ((x02 & (((x22 | x23 | (~x22 & ~x23)) & (x04 ? (x05 & ~x14) : x14)) | (x04 & x05 & x14))) | (~x14 & (x04 ? ~x02 : x05))) : ((~x02 & (~x04 | (x04 & x14))) | (x04 & x05 & ~x14) | (x02 & ~x04 & x14)))) | (x05 & ((~x14 & ((~x00 & x04 & ((x23 & ~x24 & x02 & ~x03) | (~x02 & x03 & x19 & x35))) | (~x17 & x18 & ~x20 & x02 & x03 & ~x04))) | (~x00 & ~x02 & ~x03 & x04 & x14 & x16))));
  assign z2 = x01 & ((~x05 & ((~x00 & ((~x03 & (x04 ? (x02 ? (~x14 & ((~x17 & (((~x22 | ~x23) & (~x21 | (x18 & x19 & ~x20))) | (x22 & x23 & (~x21 | (x21 & x34))) | (x21 & x34 & (~x18 | ~x19 | x20)))) | (x17 & x19 & x13 & x16))) : (x14 | (~x14 & x16))) : (x02 ? (x14 & ((x16 & (~x17 | ~x19)) | (~x16 & (x17 | x19)) | (~x17 & x19) | ~x25 | (x17 & ~x19))) : ((x06 & x07 & x09 & (~x08 | (x08 & ~x11 & (~x10 | x13)))) | (~x14 & x32))))) | (~x02 & x03 & x14 & x19 & ((x27 & x28) | (x04 & x26 & (~x22 | ~x23) & (~x27 | ~x28)))))) | (x00 & ~x02 & x03 & x14) | (~x14 & ((x00 & x02 & (~x03 | (x03 & (x22 | x23 | (~x22 & ~x23))))) | (~x02 & ((x00 & (x03 ^ x04)) | (x03 & x04 & (~x21 | (x17 & ~x20))) | (~x03 & ~x04 & ~x32 & x33 & (~x29 | ~x30 | ~x31)))))))) | (x02 & ((x05 & (x04 ? ((~x14 & (x00 ? (x03 & (x22 | x23 | (~x22 & ~x23))) : (~x03 & ((x23 & ~x24) | (x19 & x35 & (~x23 | x24)))))) | (x00 & x03 & x14)) : ((~x17 & x18 & ~x20 & x03 & ~x14) | (~x00 & ~x03 & x13 & x14 & x17 & ~x37)))) | (x00 & ~x04 & x14 & (~x03 | (x03 & (x22 | x23 | (~x22 & ~x23))))))) | (x00 & ((~x14 & (x03 ? (x04 ? ~x02 : x05) : (x04 & x05))) | (~x02 & ~x03 & (~x04 | (x04 & x14))))) | (~x00 & ~x02 & ~x03 & ~x04 & x05 & ~x14 & x38));
  assign z3 = x01 & ((~x05 & ((~x00 & ((~x03 & (x04 ? (~x14 & (x02 ? (x17 ? ~x13 : ((~x22 | ~x23) & (~x21 | (x18 & x19 & ~x20)))) : x16)) : (x02 ? (x14 & ((x16 & (~x17 | ~x19)) | (~x16 & (x17 | x19)) | (~x17 & x19) | ~x25 | (x17 & ~x19))) : ((~x14 & x32) | (x06 & x07 & (((x08 | ~x09) & (x10 ? (~x11 & ~x13) : x11)) | (~x08 & x09) | (x08 & ~x09 & ~x11))))))) | (~x02 & x03 & x14 & ((x27 & x28) ? ~x04 : (~x04 | (x04 & x19 & x26 & (~x22 | ~x23))))))) | (x00 & ~x02 & x03 & x14) | (~x14 & ((~x04 & (x02 ? ~x03 : ((x00 & x03) | (~x03 & x29 & x30 & x31 & ~x32 & x33)))) | (x03 & ((~x02 & x04 & (~x21 | (x17 & ~x20))) | (x00 & x02 & (x22 | x23 | (~x22 & ~x23))))))))) | (x02 & ((x05 & ((~x00 & (x03 ? (~x04 & ~x14 & (x17 | ~x18 | x20)) : ((x23 & ~x24 & x04 & ~x14) | (~x04 & x14 & x17 & ~x37)))) | (x03 & ((x00 & x04 & (x14 | (~x14 & (x22 | x23 | (~x22 & ~x23))))) | (~x17 & x18 & ~x20 & ~x04 & ~x14))))) | (x00 & (x03 ? (~x04 & x14 & (x22 | x23 | (~x22 & ~x23))) : (x04 ^ x14))))) | (~x00 & ~x02 & ~x03 & ~x04 & x05 & ~x14 & x38) | (x00 & ((~x02 & ((~x03 & (~x04 | (x04 & x14))) | (x04 & ~x14))) | (x03 & ~x04 & x05 & ~x14))));
  assign z4 = x01 & ((~x05 & ((~x00 & (x03 ? ((~x02 & x04 & (x14 ? ((x27 & x28) | ((~x27 | ~x28) & (~x22 | ~x23) & (~x19 | ~x26 | (x19 & x26)))) : (x21 & x34 & (~x17 | x20)))) | (~x04 & ((x02 & x36 & (~x14 | (x14 & (~x27 | ~x28)))) | (x14 & x27 & x28)))) : (x04 ? (~x14 & (x02 ? ((x13 & x17 & (x16 | (~x16 & x36))) | (~x17 & (((~x22 | ~x23) & (~x21 | (x18 & x19 & ~x20))) | (x21 & x34 & (~x18 | ~x19 | x20 | (x22 & x23)))))) : x16)) : (x02 ? (x14 & ((x16 & (~x17 | ~x19)) | (~x16 & (x17 | x19)) | (~x17 & x19) | ~x25 | (x17 & ~x19) | (x25 & (x16 ? (x17 & x19) : (~x17 & ~x19))))) : (x06 & x07 & (x08 ? (~x11 & (~x10 | (x13 & (x09 | (~x09 & x10))))) : (x09 | (~x09 & ~x10 & ~x11 & x12)))))))) | (x00 & (x02 ? (~x14 & (~x03 | (x03 & (x22 | x23)))) : (x03 ? x14 : (x04 & ~x14)))) | (~x02 & x03 & ~x04 & ~x14))) | (x02 & ((x00 & (x03 ? (((x22 | x23) & (x04 ? (x05 & ~x14) : x14)) | (x05 & (~x04 ^ x14))) : (~x04 & x14))) | (x05 & ((~x00 & ~x03 & ((x23 & ~x24 & x04 & ~x14) | (~x04 & x14 & ((x36 & x37) | (x13 & x17 & ~x37))))) | (~x17 & x18 & ~x20 & x03 & ~x04 & ~x14))))) | (~x03 & ((x04 & ((x00 & (x14 ? ~x02 : x05)) | (~x00 & ~x02 & x05 & x14 & ~x16 & x36))) | (x00 & ~x02 & ~x04))));
endmodule