module pla__in2 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18,
    z0, z1, z2, z3, z4, z5, z6, z7, z8, z9  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18;
  output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
  assign z0 = ~x00 & (x14 ? (~x15 & ((((~x07 & (x08 ? (x17 & ~x18) : (~x17 & x18))) | (x07 & ~x08 & x17 & x18)) & (~x06 ^ x16)) | (~x06 & x07 & x08 & x16 & ~x17 & ~x18))) : ((~x16 & ((~x17 & ((x10 & ((x01 & ~x11 & ~x15 & ~x18 & (~x12 | (x12 & ~x13))) | (x15 & x18))) | (~x02 & ~x06 & ~x07 & ~x10 & x15 & x18 & (~x08 | ~x09)))) | (x15 & x17 & ((~x02 & ~x06 & ~x10 & (x07 ? ((~x08 & (~x09 | x18)) | (~x09 & x18)) : (x08 & ~x18))) | (x10 & ~x18))))) | (~x02 & ~x10 & x15 & x16 & ((x08 & ~x18 & (x06 ? (~x07 & x17) : (x07 & ~x17))) | (x06 & ((~x08 & (~x09 | x18)) | (~x09 & x18)) & (~x07 ^ x17))))));
  assign z1 = x00 | (~x14 & x15 & ((~x00 & ~x02 & ~x10 & (x06 ? (x16 & ((((~x08 & (~x09 | x18)) | (~x09 & x18)) & (~x07 ^ x17)) | (x17 & ~x18 & ~x07 & x08))) : ((x08 & ~x18 & (x07 ? (x16 & ~x17) : (~x16 & x17))) | (~x16 & ((x18 & (~x08 | ~x09) & (~x07 ^ x17)) | (x07 & ~x08 & ~x09 & x17)))))) | (~x16 & ~x17 & ~x18)));
  assign z2 = ~x00 & ~x14 & ~x15 & ((((~x07 & (x08 ? (x17 & ~x18) : (~x17 & x18))) | (x07 & ~x08 & x17 & x18)) & (~x06 ^ x16) & (x09 ? x03 : x04)) | (x03 & ((~x09 & (((~x08 ^ x18) & ((x06 & x16 & (~x07 ^ x17)) | (~x16 & x17 & ~x06 & x07))) | (~x06 & ~x07 & x08 & ~x16 & ~x17 & x18))) | (~x06 & x07 & x08 & ~x17 & ~x18 & x09 & x16))) | (~x17 & ~x18 & ((x04 & ~x06 & x07 & x08 & ~x09 & x16) | (x01 & ~x03 & ~x10 & ~x16))));
  assign z3 = ~x00 & ~x14 & ~x15 & ((x03 & ((x16 & (x18 | (~x17 & ~x18))) | (x01 & x05 & ~x10) | x17 | (~x16 & ~x17 & x18))) | (x01 & ~x10 & ~x16 & ~x17 & ~x18 & (x02 | (x04 & ~x05))));
  assign z4 = ~x00 & ~x16 & ~x17 & ((x18 & ((~x15 & ((x04 & ~x06 & ~x07 & (x08 ? ~x09 : ~x14)) | (x14 & (x06 | x07 | x08)) | (x03 & ~x14))) | (~x14 & x15 & (x02 | x06 | x07 | x10 | (x08 & x09))))) | (x01 & ~x11 & ~x12 & ~x14 & ~x15 & ~x18 & (~x03 | x05 | x10)));
  assign z5 = ~x00 & ~x15 & ((~x17 & ((x07 & ((x14 & x18) | (x04 & ~x06 & x08 & x09 & ~x14 & x16 & ~x18))) | (~x07 & ((x04 & ((x18 & (~x06 ^ x16) & (x08 ? ~x09 : (x09 & ~x14))) | (x06 & ~x08 & ~x09 & x16 & ~x18))) | (x14 & x16 & ~x18))) | (x14 & ((x06 & (~x16 ^ ~x18)) | (x08 & ~x16 & x18) | (~x08 & x16 & ~x18))) | (x01 & x03 & ~x05 & ~x10 & ~x14 & ~x16 & ~x18 & ((x11 & (~x13 | (~x12 & x13))) | (x12 & (~x13 | (~x11 & x13))))))) | (x17 & ((x04 & (~x06 ^ x16) & ((x08 & ((x07 & ~x09 & x18) | (~x07 & x09 & ~x14 & ~x18))) | (x07 & ~x08 & (x09 ? (~x14 & x18) : ~x18)))) | (x14 & ((x18 & (~x07 | x08)) | (~x18 & (x07 | ~x08 | (~x06 & x16))) | (x06 & ~x16))))) | (x14 & x16 & x18 & (~x06 | x08)));
  assign z6 = ~x00 & ~x14 & ((~x17 & (((~x16 ^ ~x18) & (x15 ? (x02 | x10) : x03)) | (x15 & ((x06 & ((~x16 & x18) | (x07 & x16 & ~x18))) | (x08 & ((x09 & ~x16 & x18) | (~x07 & x16 & ~x18))) | (~x08 & x16 & ~x18 & (~x06 | x09)) | (x07 & x18))) | (~x15 & ((x04 & ~x09 & ((~x06 & ((~x07 & ~x08 & ~x16 & x18) | (x07 & x08 & x16 & ~x18))) | (x06 & ~x07 & ~x08 & x16 & x18))) | (x01 & ~x16 & ~x18 & ((~x03 & ((x11 & (~x13 | (~x12 & x13))) | (x12 & ~x13) | (~x11 & (~x12 | (x12 & x13))))) | ((x05 | x10) & (~x11 | (x11 & (~x13 | (~x12 & x13))))))))))) | ((x15 ? (x02 | x10) : x03) & (x17 | (x16 & x18))) | (x17 & ((x15 & ((~x07 & (x18 | (~x08 & ~x18))) | (x08 & (x18 ? x09 : x07)) | (x06 & ~x16) | (~x18 & ((~x06 & x16) | (~x08 & x09))))) | (x04 & ~x09 & ~x15 & (~x06 ^ x16) & (x07 ? (~x08 & x18) : (x08 & ~x18))))) | (x15 & x16 & x18 & (~x06 | (x08 & x09))));
  assign z7 = ~x00 & ((~x14 & (x15 ? (x16 & ((~x06 & (x18 | (~x02 & x07 & x08 & ~x10 & ~x17 & ~x18))) | (~x17 & ((x07 & x18) | (~x02 & x06 & ~x07 & ~x10 & ((~x08 & (~x09 | x18)) | (~x09 & x18))))) | x17 | (x18 & (x02 | x10 | (x08 & x09))))) : ((x03 & ((x16 & x18) | (x01 & ~x05 & ~x10 & x11 & ~x16 & ~x17 & ~x18 & ~x12 & x13))) | (x04 & x06 & x16 & ((~x07 & (x08 ? (x17 & ~x18) : (~x17 & x18))) | (x07 & ~x08 & x17 & x18))) | (x01 & x11 & ~x16 & ~x17 & ~x18 & (x12 ? ~x13 : (x13 & (~x03 | x05 | x10))))))) | (~x15 & x16 & ((x14 & ((~x06 & (x18 | (x07 & x08 & ~x17 & ~x18))) | x17 | (x18 & (x08 | (~x17 & (x07 | (x06 & ~x07 & ~x08))))))) | (x04 & x06 & ~x09 & ((x07 & x17 & (~x08 ^ x18)) | (~x17 & x18 & ~x07 & x08))) | (x03 & x17))));
  assign z8 = ~x00 & ((~x14 & ((~x18 & (x15 ? ((~x07 & x08 & ((x16 & ~x17) | (~x02 & ~x10 & x17 & (~x06 ^ x16)))) | (x16 & ~x17 & ((~x08 & (~x06 | x09)) | x02 | x10 | (x06 & x07)))) : (~x17 & ((x01 & ~x16 & (x11 ? ~x13 : (x12 & x13)) & (~x03 | x05 | x10 | (x03 & ~x05 & ~x10))) | (x16 & (x03 | (x07 & x08 & x04 & ~x06))))))) | (x17 & ((x07 & ~x08 & (~x06 ^ x16) & ((~x02 & ~x09 & ~x10 & x15) | (x04 & ~x15 & x18))) | (x18 & (x15 | (x03 & ~x15))))))) | (~x15 & ((x17 & ((x14 & x18) | (x08 & (~x06 ^ x16) & ((~x09 & x18 & x04 & x07) | (~x07 & x14 & ~x18))))) | (x16 & ~x17 & ~x18 & ((x06 & (x14 | (x04 & ~x07 & ~x08 & ~x09))) | (x14 & (~x07 | ~x08)))))));
  assign z9 = ~x00 & (x18 ? ((~x07 ^ x17) & (~x06 ^ x16) & ((~x02 & ~x10 & ~x14 & x15 & (~x08 | ~x09)) | (~x08 & x14 & ~x15))) : (((x17 | (x16 & ~x17)) & ((~x08 & ((x09 & ~x14 & x15) | (x14 & ~x15))) | (~x14 & (x15 ? (x02 | x10) : x03)))) | (~x15 & (x17 ? ((x04 & (~x06 ^ x16) & (x07 ? (~x08 & ~x09) : (x08 & ~x14))) | (x14 & (x07 | (~x06 & x16) | (x06 & ~x16)))) : ((~x14 & ((x01 & ~x13 & ~x16 & (((x11 | x12) & (~x03 | (x03 & ~x05 & ~x10))) | ((x05 | x10) & (x11 | (~x11 & x12))))) | (x04 & ~x06 & x07 & x08 & x16))) | (x16 & ((x06 & (x14 | (x04 & ~x07 & ~x08 & ~x09))) | (~x07 & x14)))))) | (~x14 & x15 & ((x06 & ((~x16 & x17) | (x07 & x16 & ~x17))) | (x16 & ((~x06 & (x17 | (~x08 & ~x17))) | (~x07 & x08 & ~x17))) | (x17 & (~x07 ^ x08))))));
endmodule