module pla__lin_rom ( 
    x0, x1, x2, x3, x4, x5, x6,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35  );
  input  x0, x1, x2, x3, x4, x5, x6;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35;
  assign z00 = (x6 & ((x1 & ((~x3 & ((x0 & x2 & ~x4 & x5) | (~x0 & ~x2 & ~x5))) | (~x0 & ((~x4 & x5 & ~x2 & x3) | (x2 & x4 & ~x5))) | (x0 & ((x4 & (x2 ? x3 : (~x5 | (x3 & x5)))) | (x3 & ~x4 & ~x5))))) | (~x1 & ((~x2 & ((x3 & ~x4 & ~x5) | (x0 & x5))) | (x2 & ((x4 & (x0 ? (~x3 ^ x5) : (x3 & ~x5))) | (~x0 & ~x4 & (~x3 | (x3 & x5))))) | (~x4 & ~x5 & x0 & ~x3))) | (~x0 & x2 & ~x3 & x4 & x5))) | (~x6 & ((x0 & ((~x4 & ((x1 & (x2 ? ~x5 : x3)) | (~x3 & (x5 ? ~x1 : ~x2)))) | (~x1 & x2 & x3 & x4))) | (x1 & ((~x3 & x4 & x5) | (~x0 & (x3 ? (x4 | (~x4 & x5)) : ~x4)))) | (x4 & ~x5 & ~x1 & ~x3))) | (x3 & ((~x1 & ~x5 & ((~x2 & x4) | (~x0 & x2 & ~x4))) | (x0 & x1 & x2 & ~x4 & x5)));
  assign z01 = (~x2 & ((~x0 & ((~x3 & ~x4 & x6) | (x1 & x3 & x4 & ~x5 & ~x6))) | (x6 & ((x0 & (x5 ? (x3 ? (~x4 | (~x1 & x4)) : x4) : (x1 ? (~x4 | (x3 & x4)) : x4))) | (~x4 & ~x5 & ~x1 & x3))) | (~x1 & ~x6 & ((x4 & (~x5 | (x3 & x5))) | (~x3 & x5))))) | (x2 & ((x0 & (x6 ? (x1 ? (x3 ? ~x4 : x5) : (x3 ? (x4 ^ x5) : (x4 ^ ~x5))) : ((~x3 & ~x4 & x5) | (x1 & x4 & ~x5)))) | (~x1 & ((~x0 & ((x6 & (x3 ? (x4 ^ ~x5) : (x4 ^ x5))) | (x3 & x5 & ~x6))) | (~x6 & (x3 ? (~x4 & ~x5) : (x4 & x5))))) | (~x0 & x1 & (x3 ? (x4 ? x6 : ~x5) : (x5 ? ~x4 : x6))))) | (x0 & x1 & x3 & ~x6 & (~x4 | (x4 & x5)));
  assign z02 = (x6 & ((x0 & ((~x1 & ((~x4 & x5 & ~x2 & x3) | (~x3 & x4 & ~x5))) | (x1 & (x2 ? (x5 & (~x3 ^ x4)) : (x3 & ~x5))) | (~x2 & ~x3 & x5))) | (~x0 & ((x3 & (x1 ? (x2 & ~x5) : (x4 ? ~x2 : ~x5))) | (x2 & ~x4 & x5) | (x1 & ~x3 & x4 & (x2 ^ ~x5)))) | (~x4 & ~x5 & ~x1 & ~x3) | (x1 & ~x2 & x3 & x4 & x5))) | (~x6 & (x1 ? ((~x2 & ~x5 & ((x3 & ~x4) | (x0 & ~x3 & x4))) | (~x0 & (x3 ? x5 : (~x4 | (x4 & x5))))) : ((x4 & ((x0 & (x5 ? ~x3 : x2)) | (~x5 & ((~x2 & x3) | (~x0 & (~x3 | (x2 & x3))))))) | (x0 & (x2 ? (~x4 & x5) : (x3 ? x5 : ~x4)))))) | (x0 & x2 & ((x4 & x5 & ~x1 & x3) | (x1 & ~x4 & ~x5)));
  assign z03 = (~x1 & ((x2 & (x5 ? ((x0 & (x6 | (x3 & ~x6))) | (~x0 & ~x3 & ~x4 & ~x6)) : ((x4 & (~x6 | (~x3 & x6))) | (~x0 & x3 & x6)))) | (~x3 & ((~x2 & ~x4 & x6) | (x5 & ~x6 & x0 & x4))) | (x3 & ((x0 & ((~x2 & x4 & (x5 | (~x5 & x6))) | (~x4 & ~x5 & x6))) | (~x2 & ~x4 & ~x6))))) | (x6 & (x0 ? (((x3 ^ x4) & (x2 ? x1 : x5)) | (x1 & (x3 ? (x4 & x5) : ~x4))) : (~x5 & ((x2 & ((~x3 & ~x4) | (x1 & x3 & x4))) | (x1 & ~x2 & (x3 | (~x3 & x4))))))) | (~x6 & ((x1 & ((~x0 & ((x2 & ((x4 & ~x5) | (x3 & ~x4 & x5))) | (x4 & x5 & (~x3 | (~x2 & x3))))) | (~x2 & ((~x3 & (x4 ^ x5)) | (x4 & ~x5 & x0 & x3))))) | (~x3 & ~x4 & ~x5)));
  assign z04 = (~x0 & ((~x3 & (x4 ? ((~x1 & (x2 ? x6 : x5)) | (x2 & ~x5 & ~x6)) : ((x2 & x5 & x6) | (~x5 & ~x6 & x1 & ~x2)))) | (x2 & ((x1 & ((x5 & ~x6) | (x3 & (x6 ? x4 : ~x5)))) | (~x4 & ~x5 & (x6 | (~x1 & ~x6))))) | (~x2 & ((x6 & ((x1 & (x5 ? x3 : x4)) | (x4 & ~x5 & ~x1 & x3))) | (~x1 & x3 & x5 & ~x6))))) | (x0 & ((x1 & (x2 ? ((x6 & (x3 ? (x4 ^ ~x5) : (x4 | (~x4 & x5)))) | (~x4 & ~x5 & ~x6)) : ((~x3 & (x4 ? x5 : x6)) | (x3 & x4) | (~x4 & x5 & ~x6)))) | (~x1 & (x3 ? (x2 ? (x4 ? (~x5 & x6) : x5) : (~x5 & (~x6 | (~x4 & x6)))) : (x4 & (x5 ? (x2 ^ x6) : x6)))) | (x4 & ~x5 & ~x6 & ~x2 & ~x3))) | (~x1 & ~x2 & ~x3 & ~x4 & (x5 | (~x5 & x6)));
  assign z05 = (x6 & ((x0 & (x1 ? ((x3 & x4) | (~x4 & x5 & ~x2 & ~x3)) : (x2 & (x3 ? (~x4 & x5) : ~x5)))) | (~x5 & ((x1 & ((~x0 & x2 & ~x3) | (~x2 & x3 & ~x4))) | (~x3 & x4 & ~x1 & ~x2))) | (~x1 & (x3 ? ((~x2 & x5) | (~x0 & x2 & (~x4 | (x4 & x5)))) : ((~x0 & ~x4) | (x2 & x4 & x5)))))) | (x1 & ((~x0 & x3 & (x2 ? (x5 & ~x6) : (x4 & ~x5))) | (~x3 & ~x6 & (x4 ? (~x5 | (x2 & x5)) : x5)))) | (~x1 & ((~x3 & (x2 ? (~x6 & (x4 ^ x5)) : (x4 & x5))) | (~x2 & x3 & x4 & ~x6))) | (x0 & x2 & x3 & x5 & ~x6);
  assign z06 = (x6 & (((~x2 ^ x4) & (x0 ? (~x1 & ~x3) : (x1 & ~x5))) | (~x2 & ((~x0 & ((~x3 & (x5 ? x1 : x4)) | (~x1 & x3 & x5))) | (x4 & ~x5 & ~x1 & x3) | (x0 & ((x4 & x5 & ~x1 & x3) | (x1 & (x5 ? x3 : x4)))))) | (x2 & ((x3 & (x0 ? (~x5 & (~x1 ^ x4)) : (x1 ? (~x4 & x5) : x4))) | (~x4 & ((~x1 & (x5 ? ~x3 : ~x0)) | (x0 & x1 & ~x5))))))) | (x0 & (x1 ? ((x2 & ((x3 & (x5 ? x4 : ~x6)) | (~x4 & x5) | (~x3 & x4 & ~x6))) | (~x3 & ~x4 & ~x5 & ~x6)) : ((~x2 & (x4 ? (x3 ? ~x6 : x5) : (x5 & ~x6))) | (x2 & ~x4 & ~x5 & ~x6)))) | (~x0 & ~x6 & (x2 ? (x5 | (~x1 & x4 & ~x5)) : (~x5 & (~x4 | (x1 & x4)))));
  assign z07 = x6 ? (x1 ? ((~x2 & ((~x3 & x4 & ~x5) | (~x0 & x3 & x5))) | (~x0 & (~x4 | (x4 & x5)) & (~x3 | (x2 & x3))) | (x0 & x2 & ~x3 & ~x5)) : ((~x2 & ((~x3 & ~x4) | (x0 & x3 & x5))) | (~x0 & x3 & ~x5) | (x0 & ((~x3 & x4 & x5) | (x2 & ((~x4 & x5) | (x3 & (~x5 | (x4 & x5))))))))) : ((x4 & ((x0 & ((~x2 & x5) | (x1 & x3 & ~x5))) | (~x0 & ((x1 & (x2 ? (x3 & ~x5) : x5)) | (~x1 & x2 & ~x3 & x5))) | (~x1 & ~x5 & (~x2 ^ x3)))) | (~x4 & ~x5) | (x5 & ((~x1 & ((~x2 & ~x4) | (~x0 & x2 & x3))) | (x3 & ~x4 & x1 & ~x2))));
  assign z08 = (x2 & ((x0 & ((x1 & ((~x3 & (x4 ? ~x6 : x5)) | (~x5 & x6 & (~x4 | (x3 & x4))))) | (~x1 & (x3 ? (x6 ? ~x4 : x5) : (x6 & (x4 ^ x5)))) | (~x5 & ~x6 & x3 & ~x4))) | (~x1 & ((x3 & ((x4 & ~x5 & ~x6) | (x5 & x6 & ~x0 & ~x4))) | (~x0 & ~x3 & (~x5 | (x4 & x5 & x6))))) | (~x0 & x1 & ((x3 & (~x6 | (~x4 & ~x5 & x6))) | (~x3 & ~x4 & x5 & x6))))) | (~x2 & ((x1 & ((x4 & ((~x0 & (~x3 ^ x6)) | (x6 & (x5 ? ~x3 : x0)))) | (x0 & (x3 ? (x5 & x6) : (~x5 & ~x6))) | (~x3 & ~x4 & (~x5 ^ ~x6)))) | (x4 & ((x0 & ((~x1 & x3 & x6) | (~x3 & x5 & ~x6))) | (x3 & x5 & x6 & ~x0 & ~x1))) | (~x1 & ((~x3 & ~x4 & x5 & x6) | (x3 & ~x5 & (~x6 | (~x4 & x6))))))) | (x3 & x5 & ~x6 & ~x0 & ~x1);
  assign z09 = (x6 & ((x1 & ((x0 & ((~x2 & x3 & x5) | (x4 & ~x5 & x2 & ~x3))) | (~x3 & ((~x2 & x4 & x5) | (~x0 & ~x4 & ~x5))) | (~x2 & ((~x0 & x5 & (~x4 | (x3 & x4))) | (x3 & x4 & ~x5))) | (x3 & ~x4 & ~x5 & ~x0 & x2))) | (~x1 & (x2 ? ((~x3 & ~x4 & ~x5) | (x5 & (x0 ? (x3 & ~x4) : (~x4 | (x3 & x4))))) : (x4 & ~x5))) | (x0 & ~x4 & (x2 ? (x3 & ~x5) : ~x3)))) | (x4 & ((x5 & (x1 ? (~x3 & ~x6) : (x2 ? ~x3 : (x3 & ~x6)))) | (x3 & ~x5 & ~x6 & (x1 ? (x0 | (~x0 & x2)) : x2)))) | (~x3 & ~x4 & x5 & ~x6);
  assign z10 = (x1 & ((~x5 & ((~x0 & x2 & ~x3) | (~x2 & x3 & ~x4))) | (~x0 & ((~x2 & ((~x4 & x5 & x6) | (x3 & x4 & ~x6))) | (x5 & ((x2 & (x3 ? (x4 | (~x4 & x6)) : (x4 & x6))) | (x3 & ~x4 & ~x6))))) | (x0 & ((x2 & (x3 ? (~x6 | (~x4 & x6)) : (x6 & (x4 | (~x4 & x5))))) | (~x2 & x3 & x4 & x6))))) | (~x2 & ((~x1 & ((~x3 & ((~x5 & ~x6) | (x4 & (x5 ? ~x0 : x6)))) | (x3 & ~x4 & x5 & x6))) | (x0 & ((~x3 & ~x4 & x5 & x6) | (x3 & ~x6 & (x4 | (~x4 & x5))))))) | (~x1 & ((x2 & ((x4 & ((~x0 & (x3 ? (x5 & x6) : ~x6)) | (x6 & (x5 ? x0 : x3)))) | (x0 & ~x3 & (~x6 | (~x5 & x6))) | (~x4 & ~x5 & ~x6 & ~x0 & x3))) | (~x0 & ~x3 & ~x4 & (~x5 ^ ~x6))));
  assign z11 = (x4 & (((x2 ? x6 : (x3 & ~x6)) & (x1 ? ~x0 : ~x5)) | (x6 & ((x1 & ((x0 & x2 & x3) | (~x2 & ~x3 & ~x5))) | (x0 & x2 & x5 & (~x3 | (~x1 & x3))))) | (~x3 & ~x5 & ~x6) | (x5 & (x2 ? (x3 & ~x6) : (x0 ? (x3 & ~x6) : (~x1 & ~x3)))))) | (x6 & ((x5 & (x0 ? (x2 & ~x4) : (x1 ? (x2 & ~x4) : (~x2 & x3)))) | (~x4 & ~x5 & ((~x2 & x3) | (x1 & x2 & ~x3))))) | (~x4 & ~x6 & (~x5 | (x3 & x5)));
  assign z12 = (x5 & (x4 ? ((x3 & ((~x2 & ((x0 & (~x6 | (x1 & x6))) | (~x0 & x1) | (~x1 & x6))) | (x2 & ~x6 & ~x0 & ~x1))) | (x2 & ~x3 & x6 & (x0 | (~x0 & x1)))) : ((x0 & ((~x2 & x3 & x6) | (x1 & x2 & ~x6))) | (~x2 & ((~x0 & x3 & (~x1 | (x1 & x6))) | (~x1 & ~x3 & x6))) | (~x1 & x2 & (~x3 ^ x6))))) | (x2 & ((x0 & ((~x3 & ~x4 & ~x5) | (~x1 & x3 & x4 & ~x6))) | (x4 & ((~x0 & ~x6 & (x1 ? x3 : ~x5)) | (~x5 & x6 & (~x1 | (x1 & x3))))) | (~x0 & x1 & ~x3 & ~x4 & (~x6 | (~x5 & x6))))) | (~x2 & ((~x3 & x4 & ~x6) | (~x5 & (x3 ? (x1 ? (x4 & ~x6) : ~x4) : (x4 & x6)))));
  assign z13 = (x6 & (x2 ? (x1 ? ((x0 & (x4 ? x3 : ~x5)) | (x3 & ((~x4 & x5) | (~x0 & (~x5 | (x4 & x5)))))) : (x5 ? (x0 ? x4 : ~x3) : x3)) : (x3 ? (~x4 & ~x5) : (x4 ? (~x1 | (x1 & x5)) : x5)))) | (x5 & ~x6 & (x3 ? (~x4 | (~x1 & ~x2 & x4)) : x4));
  assign z14 = (x3 & ((x1 & (x4 ? (x0 ? (x6 ? x5 : x2) : (x2 ? x5 : (~x5 & x6))) : ((~x0 & (x2 ? ~x5 : (x5 & ~x6))) | (~x2 & ~x5) | (x2 & x5 & x6)))) | (~x1 & (x2 ? ((x0 & (x4 ? (x5 & x6) : ~x6)) | (~x4 & ((~x5 & x6) | (~x0 & x5 & ~x6)))) : (x4 & (x6 ? ~x5 : ~x0)))) | (~x4 & x5 & ~x6 & x0 & ~x2))) | (~x3 & (x6 ? ((x0 & (x2 ? (x4 & ~x5) : (~x4 & x5))) | (~x0 & x1 & ((~x4 & x5) | (x2 & x4 & ~x5))) | (~x2 & (x4 ^ ~x5)) | (~x4 & x5 & ~x1 & x2)) : (~x2 ^ x4))) | (~x0 & ~x1 & x2 & (x4 ? (x5 & x6) : (~x5 & ~x6)));
  assign z15 = (x5 & (x3 ? ((x4 & ~x6 & ((x0 & (~x2 | (x1 & x2))) | (~x1 & x2) | (~x0 & x1))) | (x6 & ((~x2 & ~x4) | (~x0 & ~x1 & x2)))) : ((~x4 & ~x6) | (x2 & x6 & (x0 | (~x0 & x1)))))) | (~x5 & ~x6) | (x6 & ((~x2 & (x3 ? x4 : (~x4 & ~x5))) | (~x3 & ~x5 & (x1 ? x4 : x2))));
  assign z16 = (x4 & (x2 ? ((~x6 & (x0 ? ((~x3 & x5) | (x1 & x3 & ~x5)) : (x1 ? x5 : ~x3))) | (~x1 & (x3 ? x5 : (~x5 & x6))) | (x1 & x3 & x5 & x6)) : (x3 ? (x5 & ~x6 & (x0 | (~x0 & x1))) : ~x5))) | (~x4 & ((x1 & (x3 ? ~x5 : (x5 & x6))) | (~x1 & x2 & (x5 ? x6 : x3)) | (x5 & ((~x3 & ~x6) | (~x2 & x3 & x6))))) | (x3 & x5 & ~x6 & ~x0 & ~x1 & ~x2);
  assign z17 = (x5 & ((x6 & (x2 ? ((~x4 & ((x0 & (~x3 | (x1 & x3))) | (~x1 & x3) | (~x0 & x1))) | (~x1 & ~x3 & x4)) : ((x3 & ~x4) | (x1 & ~x3 & x4)))) | (x3 & x4 & ~x6 & (x1 | (~x1 & x2))))) | (x6 & ((~x4 & ~x5) | (~x3 & x4 & ~x1 & ~x2)));
  assign z18 = (x5 & ((x1 & ((x2 & ((x0 & (x3 ? ~x6 : (x4 & x6))) | (x3 & ~x4 & x6))) | (~x0 & (x3 ? ((~x4 & ~x6) | (~x2 & x4 & x6)) : (x4 & x6))))) | ((x3 ? (~x4 & ~x6) : (x4 & x6)) & (x2 ? ~x1 : x0)) | (~x2 & ((~x3 & x4 & ~x6) | (~x1 & x6 & (x3 ? x4 : ~x0)))))) | (~x5 & ((x4 & ((x2 & ((x6 & (x0 ? (~x3 | (x1 & x3)) : x1)) | (~x1 & x3) | (~x3 & ~x6))) | (x1 & ~x2 & x3))) | (~x3 & ~x4) | (~x1 & ~x2 & x3))) | (x3 & x4 & ~x6 & ~x0 & x1 & x2);
  assign z19 = (x4 & ((x6 & (x5 ? ((x1 & (x0 ? (x2 & x3) : (x2 | (~x2 & x3)))) | (x0 & (x2 ^ x3)) | (~x1 & x2 & x3)) : ((x1 & (~x3 | (x2 & x3))) | (~x2 & x3) | (~x1 & x2)))) | (x5 & ((~x3 & ~x6) | (~x2 & x3 & ~x0 & ~x1))))) | (~x5 & ~x6) | (~x4 & x5 & (~x6 | (~x3 & x6 & (~x2 | (~x0 & ~x1 & x2)))));
  assign z20 = (x4 & (x2 ? (x6 ? (x1 ? (~x3 & x5) : (~x3 | (x3 & x5))) : ((x0 & (x3 ? x1 : ~x5)) | (~x5 & (x1 ? ~x0 : x3)))) : (x3 ? (x5 ^ ~x6) : x6))) | (~x4 & ~x5 & x6) | (x5 & (x3 ? ((x1 & x2 & x6) | (~x2 & ~x4 & ~x6 & ~x0 & ~x1)) : (~x4 & ~x6)));
  assign z21 = x6 & (x4 ? ((~x5 & ((x1 & (~x3 | (x2 & x3))) | (~x2 & x3) | (~x1 & x2))) | (~x3 & x5 & (~x2 | (~x1 & x2)))) : x5);
  assign z22 = (x1 & ((x2 & ((x0 & x3 & (x4 ? (~x5 & x6) : (x5 & ~x6))) | (~x5 & x6 & ~x0 & x4))) | (~x4 & x5 & ~x6 & ~x0 & x3))) | (x0 & ((x4 & ~x5 & x6 & x2 & ~x3) | (~x2 & x3 & ~x4 & x5 & ~x6))) | (x3 & ((x6 & (x4 ^ x5) & (~x2 | (~x1 & x2))) | (x5 & ~x6 & (x2 ? ~x1 : x4)))) | (~x4 & ~x5 & ~x6) | (~x3 & (x4 ? (~x6 & (~x2 | (x2 & x5))) : (x5 & x6)));
  assign z23 = ~x6 | (x6 & (x4 ? ((x5 & (x2 ? ((x0 & (~x3 | (x1 & x3))) | (~x1 & x3) | (~x0 & x1)) : x3)) | (~x3 & ~x5 & ~x1 & ~x2)) : ~x5));
  assign z24 = x5 ? (~x6 & (x3 ? ((x0 & (x2 ? x1 : ~x4)) | (~x1 & x2) | (~x2 & x4) | (~x0 & x1 & (~x4 | (x2 & x4)))) : x4)) : (x6 & (~x4 | (~x3 & x4 & (~x2 | (~x1 & x2)))));
  assign z25 = x4 & x5 & x6 & (x2 ? (x1 | (~x1 & x3)) : x3);
  assign z26 = (x6 & ((x3 & ((x5 & ((~x4 & ((x0 & (~x2 | (x1 & x2))) | (~x1 & x2) | (~x0 & x1))) | (x2 & x4 & ~x0 & x1))) | (x4 & (~x2 | (x2 & (~x1 | (x0 & x1))))))) | (x4 & ((~x3 & x5) | (x2 & ~x5 & (x0 ? ~x3 : x1)))))) | (~x5 & ~x6) | (~x4 & x5 & (~x3 | (~x2 & x3 & ~x0 & ~x1)));
  assign z27 = ~x6 | (x6 & (~x5 | (x5 & (~x4 | (~x3 & x4 & (~x2 | (~x0 & ~x1 & x2)))))));
  assign z28 = x6 & (x4 ? ((x2 & (x1 ? (~x5 | (x3 & x5)) : x3)) | (~x2 & x3) | (~x3 & x5)) : x5);
  assign z30 = ~x6 | (~x5 & x6 & (~x4 | (~x3 & x4 & (~x2 | (~x0 & ~x1 & x2)))));
  assign z31 = 1'b1;
  assign z32 = 1'b1;
  assign z35 = 1'b1;
  assign z29 = 1'b0;
  assign z33 = 1'b0;
  assign z34 = 1'b0;
endmodule