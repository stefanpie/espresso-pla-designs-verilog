module pla__newxcpla1 ( 
    CPIPE1s__larrow__0__rarrow__, CPIPE1s__larrow__1__rarrow__,
    CPIPE1s__larrow__2__rarrow__, CPIPE1s__larrow__3__rarrow__,
    CPIPE1s__larrow__4__rarrow__, CPIPE1s__larrow__5__rarrow__,
    CPIPE1s__larrow__7__rarrow__, CPIPE1s__larrow__8__rarrow__, RESET,
    selaluSUM, aluCINbar1, aluselSR, selaluAND, selaluOR, selaluXOR,
    selBIbar, storeSXT, pbusLtoINB, RD_WR, predecodeEA, pSTOREwrite,
    pLOADLtobusL, pSXTtobusL, byteEX, o16, o17, o18, o19, o20, o21, o22,
    o23  );
  input  CPIPE1s__larrow__0__rarrow__, CPIPE1s__larrow__1__rarrow__,
    CPIPE1s__larrow__2__rarrow__, CPIPE1s__larrow__3__rarrow__,
    CPIPE1s__larrow__4__rarrow__, CPIPE1s__larrow__5__rarrow__,
    CPIPE1s__larrow__7__rarrow__, CPIPE1s__larrow__8__rarrow__, RESET;
  output selaluSUM, aluCINbar1, aluselSR, selaluAND, selaluOR, selaluXOR,
    selBIbar, storeSXT, pbusLtoINB, RD_WR, predecodeEA, pSTOREwrite,
    pLOADLtobusL, pSXTtobusL, byteEX, o16, o17, o18, o19, o20, o21, o22,
    o23;
  assign selaluSUM = (~CPIPE1s__larrow__4__rarrow__ & ((CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__7__rarrow__ & (CPIPE1s__larrow__3__rarrow__ | (~CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__3__rarrow__))) | (~CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__))) | (CPIPE1s__larrow__4__rarrow__ & (~CPIPE1s__larrow__3__rarrow__ | (CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__))) | ~CPIPE1s__larrow__5__rarrow__ | ~CPIPE1s__larrow__7__rarrow__ | (CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__);
  assign aluCINbar1 = CPIPE1s__larrow__7__rarrow__ & ((CPIPE1s__larrow__2__rarrow__ & ((~CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | (~CPIPE1s__larrow__2__rarrow__ & (CPIPE1s__larrow__0__rarrow__ ? (~CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__4__rarrow__) : ((~CPIPE1s__larrow__1__rarrow__ & (CPIPE1s__larrow__5__rarrow__ | (CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | (~CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__5__rarrow__)))) | (CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__3__rarrow__ & (~CPIPE1s__larrow__4__rarrow__ | ~CPIPE1s__larrow__5__rarrow__)) | (~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__));
  assign aluselSR = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__2__rarrow__;
  assign selaluAND = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__1__rarrow__;
  assign selaluOR = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__1__rarrow__;
  assign selaluXOR = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__;
  assign selBIbar = CPIPE1s__larrow__7__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__1__rarrow__ & (CPIPE1s__larrow__4__rarrow__ | (~CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__))) | (CPIPE1s__larrow__4__rarrow__ & (CPIPE1s__larrow__5__rarrow__ ? (CPIPE1s__larrow__0__rarrow__ | CPIPE1s__larrow__2__rarrow__) : ~CPIPE1s__larrow__3__rarrow__)));
  assign storeSXT = CPIPE1s__larrow__7__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__2__rarrow__;
  assign pbusLtoINB = ~CPIPE1s__larrow__7__rarrow__ | (CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__8__rarrow__ & (~CPIPE1s__larrow__3__rarrow__ | ~CPIPE1s__larrow__4__rarrow__ | ~CPIPE1s__larrow__5__rarrow__));
  assign RD_WR = (~CPIPE1s__larrow__4__rarrow__ & (CPIPE1s__larrow__2__rarrow__ ? (CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__) : (CPIPE1s__larrow__3__rarrow__ ? CPIPE1s__larrow__5__rarrow__ : (CPIPE1s__larrow__7__rarrow__ & (CPIPE1s__larrow__0__rarrow__ | (~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__5__rarrow__)))))) | ~CPIPE1s__larrow__5__rarrow__ | ~CPIPE1s__larrow__7__rarrow__ | (~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__);
  assign predecodeEA = ~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__ & (CPIPE1s__larrow__2__rarrow__ | (~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__2__rarrow__));
  assign pSTOREwrite = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__;
  assign pLOADLtobusL = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__;
  assign pSXTtobusL = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__8__rarrow__ & (~CPIPE1s__larrow__3__rarrow__ | ~CPIPE1s__larrow__4__rarrow__ | ~CPIPE1s__larrow__5__rarrow__);
  assign byteEX = CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__5__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__;
  assign o16 = (CPIPE1s__larrow__4__rarrow__ & (~CPIPE1s__larrow__3__rarrow__ | (CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__))) | ~CPIPE1s__larrow__5__rarrow__ | ~CPIPE1s__larrow__7__rarrow__ | (CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__) | (~CPIPE1s__larrow__4__rarrow__ & ((~CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (CPIPE1s__larrow__7__rarrow__ & ((CPIPE1s__larrow__0__rarrow__ & (CPIPE1s__larrow__3__rarrow__ | (~CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__3__rarrow__))) | (~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & (~CPIPE1s__larrow__2__rarrow__ | (~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__2__rarrow__))) | (CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__2__rarrow__)))))));
  assign o17 = ~CPIPE1s__larrow__5__rarrow__ | ~CPIPE1s__larrow__7__rarrow__ | (~CPIPE1s__larrow__4__rarrow__ & (CPIPE1s__larrow__2__rarrow__ ? (CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__) : (CPIPE1s__larrow__3__rarrow__ ? CPIPE1s__larrow__5__rarrow__ : (CPIPE1s__larrow__7__rarrow__ & (CPIPE1s__larrow__0__rarrow__ | (~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__5__rarrow__))))));
  assign o18 = ~CPIPE1s__larrow__5__rarrow__ | ~CPIPE1s__larrow__7__rarrow__ | (~CPIPE1s__larrow__4__rarrow__ & (CPIPE1s__larrow__2__rarrow__ ? (CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__) : (CPIPE1s__larrow__3__rarrow__ ? CPIPE1s__larrow__5__rarrow__ : (CPIPE1s__larrow__7__rarrow__ & (CPIPE1s__larrow__0__rarrow__ | (~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__5__rarrow__))))));
  assign o19 = (~CPIPE1s__larrow__5__rarrow__ & ((CPIPE1s__larrow__4__rarrow__ & ((CPIPE1s__larrow__0__rarrow__ & (CPIPE1s__larrow__1__rarrow__ | ~CPIPE1s__larrow__2__rarrow__)) | (~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__7__rarrow__))) | (~CPIPE1s__larrow__3__rarrow__ & (~CPIPE1s__larrow__0__rarrow__ | CPIPE1s__larrow__1__rarrow__)))) | (~CPIPE1s__larrow__2__rarrow__ & ((CPIPE1s__larrow__5__rarrow__ & ((~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__7__rarrow__ & (~CPIPE1s__larrow__1__rarrow__ | (~CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__4__rarrow__))) | (CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__4__rarrow__))) | (CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__7__rarrow__))) | (CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__7__rarrow__ & CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__4__rarrow__) | ~CPIPE1s__larrow__7__rarrow__ | RESET;
  assign o20 = CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__7__rarrow__ & ~RESET & ((CPIPE1s__larrow__5__rarrow__ & (CPIPE1s__larrow__0__rarrow__ | CPIPE1s__larrow__2__rarrow__)) | (~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__1__rarrow__ & ~CPIPE1s__larrow__2__rarrow__));
  assign o21 = ~RESET & CPIPE1s__larrow__7__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__2__rarrow__ & ~CPIPE1s__larrow__0__rarrow__ & ~CPIPE1s__larrow__1__rarrow__;
  assign o22 = CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__7__rarrow__ & ~RESET & ((CPIPE1s__larrow__1__rarrow__ & ((~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__) | (~CPIPE1s__larrow__0__rarrow__ & CPIPE1s__larrow__2__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__5__rarrow__))) | (~CPIPE1s__larrow__3__rarrow__ & CPIPE1s__larrow__5__rarrow__ & (CPIPE1s__larrow__0__rarrow__ | CPIPE1s__larrow__2__rarrow__)));
  assign o23 = ~RESET & CPIPE1s__larrow__7__rarrow__ & ~CPIPE1s__larrow__5__rarrow__ & CPIPE1s__larrow__4__rarrow__ & CPIPE1s__larrow__3__rarrow__ & ~CPIPE1s__larrow__1__rarrow__ & CPIPE1s__larrow__2__rarrow__;
endmodule