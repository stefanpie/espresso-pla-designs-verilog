module pla__soar.pla  ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55,
    x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69,
    x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71, z72, z73, z74, z75, z76, z77, z78, z79, z80, z81, z82, z83,
    z84, z85, z86, z87, z88, z89, z90, z91, z92, z93  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54,
    x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68,
    x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71, z72, z73, z74, z75, z76, z77, z78, z79, z80, z81, z82, z83,
    z84, z85, z86, z87, z88, z89, z90, z91, z92, z93;
  assign z00 = ~x00 | (~x01 & ~x02 & ~x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11)));
  assign z01 = ~x00;
  assign z02 = x00 & ~x17 & ~x18 & ~x19 & (x16 | (x13 & ~x14 & x15));
  assign z03 = ~x19 & ~x20 & (~x00 | ~x17 | ~x18);
  assign z04 = x00 & x17 & ~x19 & ((x14 & ((~x16 & x18) | (~x13 & x15 & x16 & ~x18))) | (~x16 & x18 & (x13 | x15)));
  assign z05 = (~x18 & (((x14 | ~x15) & (~x16 | (x13 & x17))) | (~x16 & (~x13 | x17)))) | (x18 & (~x17 | (~x13 & ~x14 & ~x15))) | ~x00 | x19;
  assign z06 = ~x19 & ~x18 & x17 & x16 & ~x15 & ~x14 & x00 & ~x13;
  assign z07 = x00 & x16 & x17 & ~x19 & ((x18 & (x13 | x15)) | (~x13 & x14 & ~x15));
  assign z08 = ~x21;
  assign z09 = x21 ? (x22 ^ x23) : (~x22 ^ x23);
  assign z10 = (x24 & (x21 ^ x22)) | (x21 & x22 & (~x23 | ~x24)) | (~x21 & ~x22 & (x23 | ~x24));
  assign z11 = x21 ^ ~x22;
  assign z12 = (x24 & (x21 | x22)) | (~x21 & ~x22 & ~x24);
  assign z13 = x00 & ~x16 & x17 & x18 & ~x20 & (x13 | x14 | x15);
  assign z14 = ~x20 & (x18 | (x00 & (~x13 | x14 | ~x15 | x16 | x17)));
  assign z15 = ~x10 & x12 & ((x07 & ((x08 & ~x09 & x11) | (x09 & ~x11))) | (x11 & (~x06 | (~x07 & ~x08 & x09))));
  assign z16 = x12 & ((x08 & ((x10 & (x11 | (~x07 & x09))) | (x00 & ~x09 & x11 & ((x25 & (x01 | x02 | x03 | x04 | ~x05)) | (~x26 & x27))))) | (x11 & (((x06 | x07) & (x10 | (x00 & ~x09 & ((x25 & (x01 | x02 | x03 | x04 | ~x05)) | (~x26 & x27))))) | (x00 & ~x09 & ~x10 & ((x25 & (x01 | x02 | x03 | x04 | ~x05)) | (~x26 & x27))))) | (x00 & ((x25 & (x01 | x02 | x03 | x04 | ~x05)) | (~x26 & x27)) & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x10 & (~x08 | x09)))) | (~x06 & x09 & x10 & ~x11));
  assign z17 = ~x18 | ~x00 | ~x17;
  assign z18 = x00 & ~x06 & ~x07 & ~x08 & ~x09 & x10 & x11 & x12 & x25 & (x01 | x02 | x03 | x04 | ~x05);
  assign z19 = x27 & ~x26 & x12 & x11 & x10 & ~x09 & ~x08 & ~x07 & x00 & ~x06;
  assign z20 = ~x20 & ~x00 & ~x18;
  assign z21 = x00 & ~x20 & ((x18 & ((~x13 & (~x17 | (~x14 & ~x15))) | (~x17 & (x14 ? (x15 & ~x16) : (~x15 & x16))))) | (~x16 & ~x18 & (x17 | (~x13 & x15))));
  assign z22 = ~x17 | ~x18 | ~x00 | ~x16;
  assign z23 = x00 & x16 & x17 & ~x20 & ((x14 & (x18 | (~x13 & ~x15))) | (x15 & x18));
  assign z24 = x34 & x37 & (((x35 | (~x36 & ~x38)) & ((~x32 & x33 & ((~x28 & (~x30 | ~x31)) | (x29 & x30 & ~x31) | (~x29 & ~x30 & x31))) | (~x31 & x32 & ~x33))) | (~x29 & x32 & ~x33 & ((x30 & ((x31 & ~x35 & (x36 | x38)) | (x35 & ~x36 & ~x38))) | (~x28 & ~x30 & x31 & ~x35))));
  assign z25 = ~x44 & (x43 | (~x42 & (x41 | (~x40 & ((x31 & ((~x33 & x34 & x37 & ((~x28 & ~x29 & ~x30 & x32 & (~x47 | (~x36 & ~x48 & ~x49 & ~x50))) | (~x32 & x35))) | (~x45 & x46))) | x39 | (~x45 & x46 & (~x32 | (~x28 & ~x29 & ~x30) | x33 | ~x34)))))));
  assign z26 = ~x43 & ~x44 & ((~x33 & x34 & ~x39 & ~x40 & ((x32 & ((~x28 & ~x29 & ~x30 & x31 & x37 & (~x47 | (~x36 & ~x48 & ~x49 & ~x50))) | (~x31 & (x28 | x29 | x30)))) | (x31 & ~x32 & x35 & x37))) | x41 | x42);
  assign z27 = ~x41 & ~x42 & ~x43 & ~x44 & ((~x33 & x34 & ((x32 & ((~x28 & ~x29 & ~x30 & x31 & x37 & (~x47 | (~x36 & ~x48 & ~x49 & ~x50))) | (~x31 & (x28 | x29 | x30)))) | (x31 & ~x32 & x35 & x37))) | x39 | x40);
  assign z28 = ~x39 & ~x40 & ~x41 & ~x42 & ~x43 & ~x44 & (x45 | x46) & (((~x32 | (~x28 & ~x29 & ~x30)) & (~x31 | ~x37)) | (x32 & ((x47 & (x36 | x48 | x49 | x50) & (x31 | (~x28 & ~x29 & ~x30))) | (x31 & (x28 | x29 | x30)))) | x33 | ~x34 | (~x32 & ~x35) | (x31 & ~x37));
  assign z29 = x00 & ((x13 & (~x17 | (x16 & ~x18))) | (~x14 & ((x16 & ~x18) | (~x13 & ~x15 & x18))) | (~x17 & (x15 | ~x16 | ~x18)));
  assign z30 = x51 & (x52 ? (x53 & ~x54) : (~x53 & x54));
  assign z31 = x18 & ~x17 & ~x16 & ~x15 & x00 & ~x13;
  assign z32 = (~x10 & ((x07 & ((x09 & ~x11) | (x08 & ~x09 & x11 & x12))) | (~x07 & ((x06 & x08 & ~x09 & ~x11) | (~x08 & x09 & x11 & x12))) | (~x06 & x11 & x12))) | (~x11 & ~x12);
  assign z33 = x00 & ((~x02 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11)) & (x01 | x03)) | (x12 & x25 & (x02 | x04 | ~x05) & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x10 & (~x08 | x09 | (~x09 & x11))))));
  assign z34 = (~x10 & ((x07 & ((x09 & ~x11) | (x08 & ~x09 & x11 & x12))) | (~x07 & ((x06 & x08 & ~x09 & ~x11) | (~x08 & x09 & x11 & x12))) | (~x06 & x11 & x12))) | (~x11 & ~x12);
  assign z35 = ~x20 & ~x00 & ~x18;
  assign z36 = ~x20 & ~x18 & ~x17 & x16 & x00 & x13;
  assign z37 = ~x18 & ~x17 & x16 & x00 & x15;
  assign z38 = x57 & ~x56 & ~x55 & x18 & ~x17 & x16 & x15 & ~x14 & x00 & ~x13;
  assign z39 = x57 & x56 & ~x55 & x18 & ~x17 & x16 & x15 & ~x14 & x00 & ~x13;
  assign z40 = x57 & ~x56 & x55 & x18 & ~x17 & x16 & x15 & ~x14 & x00 & ~x13;
  assign z41 = x57 & x56 & x55 & x18 & ~x17 & x16 & x15 & ~x14 & x00 & ~x13;
  assign z42 = x57 & ~x56 & ~x55 & x18 & ~x17 & x16 & x15 & x14 & x00 & ~x13;
  assign z43 = x57 & x56 & ~x55 & x18 & ~x17 & x16 & x15 & x14 & x00 & ~x13;
  assign z44 = x57 & ~x56 & x55 & x18 & ~x17 & x16 & x15 & x14 & x00 & ~x13;
  assign z45 = x57 & x56 & x55 & x18 & ~x17 & x16 & x15 & x14 & x00 & ~x13;
  assign z46 = ~x20 & (~x00 | ~x13 | x14 | ~x15 | x16 | x17 | x18);
  assign z47 = ~x11 & (~x12 | (x06 & ~x07 & x08 & ~x09 & ~x10));
  assign z48 = x12 & ~x11 & ~x10 & x07 & x09;
  assign z49 = ~x20 & ((x15 & ((x17 & x18) | (~x14 & x16 & ~x18))) | (x16 & ~x18 & (~x13 | ~x17)) | ~x00 | (x17 & x18 & (x13 | x14)));
  assign z50 = ~x19 & ~x20 & (~x00 | (x16 & ~x17 & ~x18));
  assign z51 = (~x64 & (x60 ? ((~x59 | ~x62) & ((x51 & ((x61 & (x52 ? (x53 ? x63 : ~x54) : (x53 & ~x54))) | (~x52 & ~x53 & ~x63))) | (~x63 & (~x61 | (~x51 & ~x54))))) : ((x61 & ((~x51 & (x54 | x63)) | (x52 & ((~x53 & x54) | (x51 & x53 & ~x63))) | (~x52 & (x53 ? x54 : x63)) | (x59 & x62))) | (x59 & x62 & ~x63)))) | (x61 & ~x62 & ~x63 & (((x52 ^ x53) & ((x51 & ~x54 & ~x59 & x60) | (x54 & ~x58 & ~x60))) | (x64 & ((x60 & (x58 | (x51 & x52 & x53 & ~x59))) | (~x58 & ~x60 & (~x51 | x59 | (~x52 & ~x53)))))));
  assign z52 = ~x20 & ((~x18 & (x13 | x15)) | ~x00 | ~x16 | ~x17 | (~x15 & x18 & ~x13 & ~x14));
  assign z53 = x00 & x12 & ~x26 & x27 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x10 & (~x08 | x09 | (~x09 & x11))));
  assign z54 = x18 & x17 & x00 & x16;
  assign z55 = x12 & x11 & ~x09 & x10;
  assign z56 = x00 & ~x19 & ~x20 & ((x18 & ((~x13 & (~x17 | (~x14 & ~x15))) | (~x17 & (x14 ? (x15 & ~x16) : (~x15 & x16))))) | (~x16 & ~x18 & (x17 | (x15 & (~x13 | ~x14)))));
  assign z57 = x00 & x01 & x02 & ~x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z58 = x00 & ~x01 & x02 & ~x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z59 = x18 & x17 & x16 & ~x15 & ~x14 & x00 & ~x13;
  assign z60 = x00 & x65 & (~x16 | ~x17 | ~x18);
  assign z61 = ~x00 | (x65 & (~x16 | ~x17 | ~x18));
  assign z62 = ~x18 | ~x00 | ~x17;
  assign z63 = x00 & x02 & x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z64 = x66 | (x00 & ((x13 & ((~x15 & ((x14 & ~x17 & x18) | (x16 & x17 & ~x18))) | (x14 & ~x18 & (x16 ^ ~x17)) | (~x17 & x18 & (x16 ? x15 : ~x14)))) | (~x17 & ~x18 & ~x15 & ~x16)));
  assign z65 = ~x30 & x31 & ~x32 & x33 & x34 & x37 & (~x28 | ~x29);
  assign z66 = x00 & ~x01 & x02 & x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z67 = x00 & x01 & ~x02 & ~x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z68 = x00 & x01 & x02 & x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z69 = x00 & ~x01 & ~x02 & x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z70 = x00 & x01 & ~x02 & x03 & ~x04 & x05 & ((~x11 & (~x09 | (x06 & (x07 | ~x08)))) | ~x10 | ~x12 | (~x06 & ~x07 & ~x08 & x11));
  assign z71 = x00 & ~x14 & x16 & x17 & ~x18 & (~x13 | x15);
  assign z72 = (x70 & (((~x71 | ~x72) & (~x73 | ~x74)) | (~x71 & ~x72))) | x67 | ~x68 | x69;
  assign z73 = x12 & x75 & ~x76 & ~x77 & ~x78 & x79 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x09 & x11) | (~x10 & (~x08 | x09)));
  assign z74 = x12 & ~x75 & ~x76 & x77 & ~x78 & x79 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x09 & x11) | (~x10 & (~x08 | x09)));
  assign z75 = x12 & x75 & ~x76 & x77 & ~x78 & x79 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x09 & x11) | (~x10 & (~x08 | x09)));
  assign z76 = x00 & ((~x06 & ((x09 & x10) | (x08 & ~x09 & ~x11))) | (x08 & ((~x07 & (x09 ? x10 : ~x11)) | (x10 & x11 & x12))) | (x10 & (x11 ? (x09 | (x12 & (x06 | x07))) : ~x09)) | (~x01 & ~x02 & ~x03 & ~x04 & x05) | ~x12 | ~x25);
  assign z77 = x00 & ((~x06 & ((x09 & x10) | (x08 & ~x09 & ~x11))) | (x08 & ((~x07 & (x09 ? x10 : ~x11)) | (x10 & x11 & x12))) | (x10 & (x11 ? (x09 | (x12 & (x06 | x07))) : ~x09)) | ~x12 | x26 | ~x27);
  assign z78 = x00 & ((~x13 & x14 & (x17 | (~x15 & x16 & x18))) | (x17 & (x18 ? (x13 | x15) : ~x16)));
  assign z79 = x18 & ~x17 & ~x16 & x15 & x14 & x00 & ~x13;
  assign z80 = x18 & ~x17 & ~x16 & x15 & x14 & x00 & x13;
  assign z81 = (~x15 & (x13 | x16)) | (x13 & (~x14 | x16)) | ~x00 | x17 | ~x18;
  assign z82 = x18 & ~x17 & ~x16 & x15 & ~x14 & x00 & ~x13;
  assign z83 = x00 & ~x13 & ~x15 & ~x16 & ~x17 & x18 & ((~x80 & x81) | (x14 & x80 & x82));
  assign z84 = x00 & ~x13 & ~x15 & ~x16 & ~x17 & x18 & x81 & (x14 | x80);
  assign z85 = x34 & ~x33 & x32 & ~x31 & ~x30 & ~x28 & ~x29;
  assign z86 = ~x18 & x17 & x16 & ~x15 & x00 & ~x13;
  assign z87 = ~x18 & ~x17 & ~x16 & x15 & ~x14 & x00 & x13;
  assign z88 = (x09 & ((x06 & ~x11 & (x07 | (~x08 & x10))) | (x07 & ~x10 & x12))) | (~x11 & ~x12) | (x12 & ((x11 & (~x09 | ~x10)) | (~x09 & ~x10 & (x06 | ~x08))));
  assign z89 = x12 & ~x75 & x76 & x77 & ~x78 & x79 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x09 & x11) | (~x10 & (~x08 | x09)));
  assign z90 = x12 & x75 & x76 & x77 & ~x78 & x79 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x09 & x11) | (~x10 & (~x08 | x09)));
  assign z91 = x12 & x75 & x76 & ~x77 & ~x78 & x79 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x09 & x11) | (~x10 & (~x08 | x09)));
  assign z92 = x12 & ~x75 & x76 & ~x77 & ~x78 & x79 & ((x06 & ((x07 & (~x10 | (x09 & ~x11))) | (~x08 & x09 & ~x11))) | (~x09 & x11) | (~x10 & (~x08 | x09)));
  assign z93 = ~x19 & ~x18 & x17 & x16 & x15 & x00 & ~x14;
endmodule