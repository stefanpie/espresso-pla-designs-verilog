module pla__apla ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11;
  assign z00 = ~x0 & ~x2 & ~x3 & ((~x6 & (x1 ? (~x4 & ~x5 & (x7 ? (x8 ^ x9) : (~x8 & ~x9))) : ((~x7 & (~x9 | (x8 & x9)) & (x4 ^ x5)) | (x4 & ~x5 & x7 & ~x8 & x9)))) | (~x1 & ~x4 & ~x5 & x6 & ~x7 & x8));
  assign z01 = ~x0 & ~x2 & ~x3 & ((~x6 & (x1 ? (~x4 & ~x5 & (x7 ? (~x8 ^ x9) : (~x8 & x9))) : (x4 ? (~x5 & (x7 ? (~x9 | (x8 & x9)) : (~x8 & x9))) : (x5 & (x7 ? x8 : (~x8 & x9)))))) | (~x1 & ~x4 & ~x5 & x6 & x7 & x8));
  assign z02 = ~x4 & ~x9 & ((~x1 & ((~x5 & ((~x6 & (~x7 | (x7 & ~x8)) & (x0 ? (~x2 & ~x3) : (x2 ^ x3))) | (~x0 & ~x2 & ~x3 & x6 & ~x8))) | (~x0 & ~x2 & ~x3 & x7 & ~x8 & x5 & ~x6))) | (~x2 & ~x3 & ~x0 & x1 & ~x7 & x8 & ~x5 & ~x6));
  assign z03 = ~x1 & ~x4 & ~x5 & ~x7 & x9 & ((~x0 & (x2 ? (~x3 & ~x6) : (~x8 & (x3 ^ x6)))) | (~x3 & ~x6 & x0 & ~x2));
  assign z04 = ~x4 & ((~x1 & ((~x5 & ((~x6 & ((x7 & (x8 ^ x9) & (x0 ? (~x2 & ~x3) : (x2 ^ x3))) | (~x0 & ~x2 & x3 & ~x7 & x8 & x9))) | (~x0 & ~x2 & ~x3 & ~x8 & x9 & x6 & x7))) | (~x0 & ~x2 & ~x3 & x5 & ~x8 & x9 & ~x6 & x7))) | (~x2 & ~x3 & ~x0 & x1 & ~x5 & ~x6 & ~x7 & x8 & x9));
  assign z05 = ~x1 & ~x3 & ~x4 & ~x5 & ~x6 & x7 & x8 & x9 & (~x0 ^ ~x2);
  assign z06 = x9 & x8 & x7 & ~x6 & ~x5 & ~x4 & x3 & ~x2 & ~x0 & ~x1;
  assign z07 = ~x0 & ~x1 & ((~x4 & ((~x6 & ((~x3 & ((~x8 & (x2 ? (~x5 & (~x7 | (x7 & x9))) : (x5 & x7))) | (~x2 & x5 & x8))) | (~x2 & x3 & ~x5 & x7 & (~x9 | (x8 & x9))))) | (~x2 & ~x3 & ~x5 & x6))) | (~x2 & ~x3 & x4 & ~x5 & ~x6 & x8));
  assign z08 = ~x3 & ~x6 & ((~x1 & (x0 ? (~x2 & ~x4 & ~x5 & (x7 ? (~x9 | (x8 & x9)) : x8)) : ((~x7 & ((~x2 & ~x8 & (x4 ^ x5)) | (x2 & ~x4 & ~x5 & x8))) | (x2 & ~x4 & ~x5 & x7 & (~x9 | (x8 & x9)))))) | (~x0 & x1 & ~x2 & ~x4 & ~x5 & ~x7 & ~x8));
  assign z09 = ~x0 & ~x2 & ((~x3 & ((~x4 & ((~x5 & (x1 ? (~x6 & (x7 ^ x8)) : (x6 & ((x8 & x9) | (x7 & ~x8 & ~x9))))) | (~x1 & x5 & ~x6 & (x8 ? x9 : x7)))) | (~x1 & x4 & ~x5 & ~x6 & (x8 ? x9 : x7)))) | (~x1 & x3 & ~x4 & ~x5 & ~x6 & (x7 ? ~x9 : x8)));
  assign z10 = ~x1 & ~x4 & ~x5 & (x0 ? (~x2 & ~x3 & ~x6 & (~x7 | (x7 & (x8 ^ x9)))) : ((~x8 & ((~x2 & (x3 ^ x6) & (~x7 | (x7 & x9))) | (x2 & ~x3 & ~x6 & x7 & x9))) | (x2 & ~x3 & ~x6 & (~x7 | (x7 & x8 & ~x9)))));
  assign z11 = ~x0 & ~x2 & ~x3 & ((~x4 & ((~x6 & (x1 ? (~x5 & (~x8 | (x7 & x8))) : (x5 & (~x7 | (x7 & x8))))) | (~x1 & ~x5 & x6 & x8))) | (~x5 & ~x6 & ~x1 & x4));
endmodule