module pla__apex5 ( 
    x000, x001, x002, x003, x004, x005, x006, x007, x008, x009, x010, x011,
    x012, x013, x014, x015, x016, x017, x018, x019, x020, x021, x022, x023,
    x024, x025, x026, x027, x028, x029, x030, x031, x032, x033, x034, x035,
    x036, x037, x038, x039, x040, x041, x042, x043, x044, x045, x046, x047,
    x048, x049, x050, x051, x052, x053, x054, x055, x056, x057, x058, x059,
    x060, x061, x062, x063, x064, x065, x066, x067, x068, x069, x070, x071,
    x072, x073, x074, x075, x076, x077, x078, x079, x080, x081, x082, x083,
    x084, x085, x086, x087, x088, x089, x090, x091, x092, x093, x094, x095,
    x096, x097, x098, x099, x100, x101, x102, x103, x104, x105, x106, x107,
    x108, x109, x110, x111, x112, x113, x114, x115, x116,
    z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71, z72, z73, z74, z75, z76, z77, z78, z79, z80, z81, z82, z83,
    z84, z85, z86, z87  );
  input  x000, x001, x002, x003, x004, x005, x006, x007, x008, x009,
    x010, x011, x012, x013, x014, x015, x016, x017, x018, x019, x020, x021,
    x022, x023, x024, x025, x026, x027, x028, x029, x030, x031, x032, x033,
    x034, x035, x036, x037, x038, x039, x040, x041, x042, x043, x044, x045,
    x046, x047, x048, x049, x050, x051, x052, x053, x054, x055, x056, x057,
    x058, x059, x060, x061, x062, x063, x064, x065, x066, x067, x068, x069,
    x070, x071, x072, x073, x074, x075, x076, x077, x078, x079, x080, x081,
    x082, x083, x084, x085, x086, x087, x088, x089, x090, x091, x092, x093,
    x094, x095, x096, x097, x098, x099, x100, x101, x102, x103, x104, x105,
    x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116;
  output z00, z01, z02, z03, z04, z05, z06, z07, z08, z09, z10, z11, z12, z13,
    z14, z15, z16, z17, z18, z19, z20, z21, z22, z23, z24, z25, z26, z27,
    z28, z29, z30, z31, z32, z33, z34, z35, z36, z37, z38, z39, z40, z41,
    z42, z43, z44, z45, z46, z47, z48, z49, z50, z51, z52, z53, z54, z55,
    z56, z57, z58, z59, z60, z61, z62, z63, z64, z65, z66, z67, z68, z69,
    z70, z71, z72, z73, z74, z75, z76, z77, z78, z79, z80, z81, z82, z83,
    z84, z85, z86, z87;
  assign z00 = x092;
  assign z01 = x099 | x100 | x097 | x098 | x095 | x096 | x093 | x094;
  assign z02 = (x036 & (x000 | ~x001 | ~x004)) | (~x000 & x001 & x004 & x028);
  assign z03 = x004 & ((x000 & x001 & ~x028 & ((~x025 & ((~x027 & (x023 ? (x024 ? (~x026 & x085) : (x026 ? x069 : x093)) : (x024 ? (~x026 & x077) : (x026 & x061)))) | (~x023 & ~x024 & ~x026 & x027 & x045))) | (~x023 & ~x024 & x025 & ~x026 & ~x027 & x053))) | (x037 & (((x025 | x027) & (x023 | x024 | x026)) | (x024 & x026) | ~x000 | ~x001 | (x025 & x027) | x028 | (~x023 & ~x024 & ~x025 & ~x026 & ~x027))));
  assign z04 = x004 & ((x000 & x001 & ~x028 & ((~x025 & ((~x027 & (x023 ? (x024 ? (~x026 & x086) : (x026 ? x070 : x094)) : (x024 ? (~x026 & x078) : (x026 & x062)))) | (~x023 & ~x024 & ~x026 & x027 & x046))) | (~x023 & ~x024 & x025 & ~x026 & ~x027 & x054))) | (x038 & (((x025 | x027) & (x023 | x024 | x026)) | (x024 & x026) | ~x000 | ~x001 | (x025 & x027) | x028 | (~x023 & ~x024 & ~x025 & ~x026 & ~x027))));
  assign z05 = x004 & ((x000 & x001 & ~x028 & ((~x025 & ((~x027 & (x023 ? (x024 ? (~x026 & x087) : (x026 ? x071 : x095)) : (x024 ? (~x026 & x079) : (x026 & x063)))) | (~x023 & ~x024 & ~x026 & x027 & x047))) | (~x023 & ~x024 & x025 & ~x026 & ~x027 & x055))) | (x039 & (((x025 | x027) & (x023 | x024 | x026)) | (x024 & x026) | ~x000 | ~x001 | (x025 & x027) | x028 | (~x023 & ~x024 & ~x025 & ~x026 & ~x027))));
  assign z06 = x004 & ((x000 & x001 & ~x028 & ((~x025 & ((~x027 & (x023 ? (x024 ? (~x026 & x088) : (x026 ? x072 : x096)) : (x024 ? (~x026 & x080) : (x026 & x064)))) | (~x023 & ~x024 & ~x026 & x027 & x048))) | (~x023 & ~x024 & x025 & ~x026 & ~x027 & x056))) | (x040 & (((x025 | x027) & (x023 | x024 | x026)) | (x024 & x026) | ~x000 | ~x001 | (x025 & x027) | x028 | (~x023 & ~x024 & ~x025 & ~x026 & ~x027))));
  assign z07 = x004 & ((x000 & x001 & ~x028 & ((~x025 & ((~x027 & (x023 ? (x024 ? (~x026 & x089) : (x026 ? x073 : x097)) : (x024 ? (~x026 & x081) : (x026 & x065)))) | (~x023 & ~x024 & ~x026 & x027 & x049))) | (~x023 & ~x024 & x025 & ~x026 & ~x027 & x057))) | (x041 & (((x025 | x027) & (x023 | x024 | x026)) | (x024 & x026) | ~x000 | ~x001 | (x025 & x027) | x028 | (~x023 & ~x024 & ~x025 & ~x026 & ~x027))));
  assign z08 = x004 & ((x000 & x001 & ~x028 & ((~x025 & ((~x027 & (x023 ? (x024 ? (~x026 & x090) : (x026 ? x074 : x098)) : (x024 ? (~x026 & x082) : (x026 & x066)))) | (~x023 & ~x024 & ~x026 & x027 & x050))) | (~x023 & ~x024 & x025 & ~x026 & ~x027 & x058))) | (x042 & (((x025 | x027) & (x023 | x024 | x026)) | (x024 & x026) | ~x000 | ~x001 | (x025 & x027) | x028 | (~x023 & ~x024 & ~x025 & ~x026 & ~x027))));
  assign z09 = x004 & ((x000 & x001 & ~x025 & ~x028 & ((~x027 & (x023 ? (x024 ? (~x026 & x091) : (x026 ? x075 : x099)) : (x024 ? (~x026 & x083) : (x026 & x067)))) | (~x023 & ~x024 & ~x026 & x027 & x051))) | (x043 & ((x024 & (x026 | x027)) | (x027 & (x023 | x026)) | ~x000 | ~x001 | x025 | x028 | (~x023 & ~x024 & ~x026 & ~x027))));
  assign z10 = x004 & ((x000 & x001 & ~x025 & ~x028 & ((~x027 & (x023 ? (x024 ? (~x026 & x092) : (x026 ? x076 : x100)) : (x024 ? (~x026 & x084) : (x026 & x068)))) | (~x023 & ~x024 & ~x026 & x027 & x052))) | (x044 & ((x024 & (x026 | x027)) | (x027 & (x023 | x026)) | ~x000 | ~x001 | x025 | x028 | (~x023 & ~x024 & ~x026 & ~x027))));
  assign z11 = x004 & ((x045 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x000 & x001 & x015 & ~x023 & ~x024 & ~x025 & ~x026 & x027 & ~x028));
  assign z12 = x004 & ((x046 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x024 & ~x025 & ~x026 & x027 & ~x028 & ~x000 & x001 & x016 & ~x023));
  assign z13 = x004 & ((x047 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x024 & ~x025 & ~x026 & x027 & ~x028 & ~x000 & x001 & x017 & ~x023));
  assign z14 = x004 & ((x048 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x024 & ~x025 & ~x026 & x027 & ~x028 & ~x000 & x001 & x018 & ~x023));
  assign z15 = x004 & ((x049 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x024 & ~x025 & ~x026 & x027 & ~x028 & ~x000 & x001 & x019 & ~x023));
  assign z16 = x004 & ((x050 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x024 & ~x025 & ~x026 & x027 & ~x028 & ~x000 & x001 & x020 & ~x023));
  assign z17 = x004 & ((x051 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x024 & ~x025 & ~x026 & x027 & ~x028 & ~x000 & x001 & x021 & ~x023));
  assign z18 = x004 & ((x052 & (x000 | ~x001 | x023 | x024 | x025 | x026 | ~x027 | x028)) | (~x024 & ~x025 & ~x026 & x027 & ~x028 & ~x000 & x001 & x022 & ~x023));
  assign z19 = x087;
  assign z20 = x088;
  assign z21 = x004 & ((x053 & (x000 | ~x001 | x023 | x024 | ~x025 | x026 | x027 | x028)) | (~x000 & x001 & x015 & ~x023 & ~x024 & x025 & ~x026 & ~x027 & ~x028));
  assign z22 = x004 & ((x054 & (x000 | ~x001 | x023 | x024 | ~x025 | x026 | x027 | x028)) | (~x000 & x001 & x016 & ~x023 & ~x024 & x025 & ~x026 & ~x027 & ~x028));
  assign z23 = x004 & ((x055 & (x000 | ~x001 | x023 | x024 | ~x025 | x026 | x027 | x028)) | (~x000 & x001 & x017 & ~x023 & ~x024 & x025 & ~x026 & ~x027 & ~x028));
  assign z24 = x004 & ((x056 & (x000 | ~x001 | x023 | x024 | ~x025 | x026 | x027 | x028)) | (~x000 & x001 & x018 & ~x023 & ~x024 & x025 & ~x026 & ~x027 & ~x028));
  assign z25 = x004 & ((x057 & (x000 | ~x001 | x023 | x024 | ~x025 | x026 | x027 | x028)) | (~x000 & x001 & x019 & ~x023 & ~x024 & x025 & ~x026 & ~x027 & ~x028));
  assign z26 = x004 & ((x058 & (x000 | ~x001 | x023 | x024 | ~x025 | x026 | x027 | x028)) | (~x000 & x001 & x020 & ~x023 & ~x024 & x025 & ~x026 & ~x027 & ~x028));
  assign z27 = x004 & x035;
  assign z28 = x004 & x034;
  assign z32 = x004 & ((x061 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x101 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x015 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z33 = x004 & ((x062 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x102 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x016 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z34 = x004 & ((x063 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x103 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x017 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z35 = x004 & ((x064 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x104 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x018 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z36 = x004 & ((x065 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x105 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x019 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z37 = x004 & ((x066 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x106 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x020 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z38 = x004 & ((x067 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x107 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x021 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z39 = x004 & ((x068 & ((x000 & (~x006 | (x001 & ~x023 & ~x024 & ~x027 & ~x028 & ~x025 & x026))) | (~x006 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)))) | (x006 & x108 & (~x001 | x023 | x024 | x027 | x028 | x025 | ~x026)) | (~x000 & x001 & x022 & ~x023 & ~x024 & ~x025 & x026 & ~x027 & ~x028));
  assign z40 = x004 & ((x069 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x109 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x015 & x023));
  assign z41 = x004 & ((x070 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x110 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x016 & x023));
  assign z42 = x004 & ((x071 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x111 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x017 & x023));
  assign z43 = x004 & ((x072 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x112 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x018 & x023));
  assign z44 = x004 & ((x073 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x113 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x019 & x023));
  assign z45 = x004 & ((x074 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x114 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x020 & x023));
  assign z46 = x004 & ((x075 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x115 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x021 & x023));
  assign z47 = x004 & ((x076 & ((x000 & (~x006 | (~x027 & ~x028 & ~x025 & x026 & x001 & x023 & ~x024))) | (~x006 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)))) | (x006 & x116 & (x027 | x028 | x025 | ~x026 | ~x001 | ~x023 | x024)) | (~x024 & ~x025 & x026 & ~x027 & ~x028 & ~x000 & x001 & x022 & x023));
  assign z48 = (x077 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x015 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z49 = (x078 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x016 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z50 = (x079 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x017 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z51 = (x080 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x018 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z52 = (x081 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x019 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z53 = (x082 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x020 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z54 = (x083 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x021 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z55 = (x084 & (x000 | ~x001 | x023 | ~x024 | x025 | x026 | x027 | x028)) | ~x004 | (~x000 & x001 & x022 & ~x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025);
  assign z56 = x004 & ((x085 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x015 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z57 = x004 & ((x086 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x016 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z58 = x004 & ((x087 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x017 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z59 = x004 & ((x088 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x018 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z60 = x004 & ((x089 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x019 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z61 = x004 & ((x090 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x020 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z62 = x004 & ((x091 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x021 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z63 = x004 & ((x092 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | ~x024)) | (~x000 & x001 & x022 & x023 & ~x026 & ~x027 & ~x028 & x024 & ~x025));
  assign z64 = x004 & ((~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x029 & x030 & x031 & x032 & ~x033 & ((~x015 & x024 & (x007 ? (x023 ? ~x077 : ~x085) : (~x023 & x085))) | (x023 & ~x077 & ~x007 & x015))) | (x015 & x023 & ~x024))) | (x029 & x030 & x031 & x032 & ~x033 & ~x077 & (x007 ^ x085) & (x025 | x026 | x027 | x028 | ~x001 | (~x023 & ~x024) | (x000 & x024))) | (x093 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | x024)));
  assign z65 = x004 & ((~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x029 & x030 & x031 & x032 & ~x033 & ((~x016 & x024 & (x008 ? (x023 ? ~x078 : ~x086) : (~x023 & x086))) | (x023 & ~x078 & ~x008 & x016))) | (x016 & x023 & ~x024))) | (x029 & x030 & x031 & x032 & ~x033 & ~x078 & (x025 | x026 | x027 | x028 | ~x001 | (~x023 & ~x024) | (x000 & x024)) & (x008 ^ x086)) | (x094 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | x024)));
  assign z66 = x004 & ((x000 & (x095 | (x009 & ~x023 & x029 & x030 & x031 & x032 & ~x033 & ~x079))) | (~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x017 & x023 & ~x024) | (~x023 & x024 & x009 & ~x017 & x029 & x030 & x031 & x032 & ~x033))) | ((x095 | (x031 & x032 & ~x033 & ~x079 & x009 & x029 & x030)) & (x026 | x027 | x028 | ~x001 | x025)) | (x009 & x029 & x030 & x031 & x032 & ~x033 & ~x079 & (x023 ^ ~x024)) | (x095 & (~x023 | x024)));
  assign z67 = x004 & ((x000 & (x096 | (x029 & x030 & x010 & ~x023 & x031 & x032 & ~x033 & ~x080))) | (~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x018 & x023 & ~x024) | (x029 & x030 & x031 & x032 & ~x033 & ~x023 & x024 & x010 & ~x018))) | ((x026 | x027 | x028 | ~x001 | x025) & (x096 | (x031 & x032 & ~x033 & ~x080 & x010 & x029 & x030))) | (x010 & x029 & x030 & x031 & x032 & ~x033 & ~x080 & (x023 ^ ~x024)) | (x096 & (~x023 | x024)));
  assign z68 = x004 & ((~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x029 & x030 & x031 & x032 & ~x033 & ((~x019 & x024 & (x011 ? (x023 ? ~x081 : ~x089) : (~x023 & x089))) | (x023 & ~x081 & ~x011 & x019))) | (x019 & x023 & ~x024))) | (x029 & x030 & x031 & x032 & ~x033 & ~x081 & (x025 | x026 | x027 | x028 | ~x001 | (~x023 & ~x024) | (x000 & x024)) & (x011 ^ x089)) | (x097 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | x024)));
  assign z69 = x004 & ((~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x029 & x030 & x031 & x032 & ~x033 & ((~x020 & x024 & (x012 ? (x023 ? ~x082 : ~x090) : (~x023 & x090))) | (x023 & ~x082 & ~x012 & x020))) | (x020 & x023 & ~x024))) | (x029 & x030 & x031 & x032 & ~x033 & ~x082 & (x025 | x026 | x027 | x028 | ~x001 | (~x023 & ~x024) | (x000 & x024)) & (x012 ^ x090)) | (x098 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | x024)));
  assign z70 = x004 & ((~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x029 & x030 & x031 & x032 & ~x033 & ((~x021 & x024 & (x013 ? (x023 ? ~x083 : ~x091) : (~x023 & x091))) | (x023 & ~x083 & ~x013 & x021))) | (x021 & x023 & ~x024))) | (x029 & x030 & x031 & x032 & ~x033 & ~x083 & (x025 | x026 | x027 | x028 | ~x001 | (~x023 & ~x024) | (x000 & x024)) & (x013 ^ x091)) | (x099 & (x025 | x026 | x027 | x028 | x000 | ~x001 | ~x023 | x024)));
  assign z71 = x004 & ((x000 & (x100 | (x029 & x030 & x014 & ~x023 & x031 & x032 & ~x033 & ~x084))) | (~x000 & x001 & ~x025 & ~x026 & ~x027 & ~x028 & ((x022 & x023 & ~x024) | (x029 & x030 & x031 & x032 & ~x033 & ~x023 & x024 & x014 & ~x022))) | ((x026 | x027 | x028 | ~x001 | x025) & (x100 | (x031 & x032 & ~x033 & ~x084 & x014 & x029 & x030))) | (x014 & x029 & x030 & x031 & x032 & ~x033 & ~x084 & (x023 ^ ~x024)) | (x100 & (~x023 | x024)));
  assign z72 = x004 & ((~x006 & x101 & (~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | (x102 & x103 & x104 & x105 & x106 & x107 & x108 & x109 & x110 & x111 & x112 & x113 & x114 & x115 & x116))) | (x003 & x029 & x030 & x031 & x032 & ~x033 & (~x101 | (x006 & (~x102 | ~x103 | ~x104 | ~x105 | ~x106 | ~x107 | ~x108 | ~x109 | ~x110 | ~x111 | ~x112 | ~x113 | ~x114 | ~x115 | ~x116)))));
  assign z73 = x004 & ~x006 & ((x101 & ((x102 & x103 & x104 & x105 & x106 & x107 & x108 & x109 & x110 & x111 & x112 & x113 & x114 & x115 & x116) | (x003 & x029 & x030 & x031 & x032 & ~x033 & ~x102))) | (x102 & (~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x101)));
  assign z74 = x004 & ~x006 & ((x101 & x102 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x103) | (x103 & x104 & x105 & x106 & x107 & x108 & x109 & x113 & x114 & x115 & x116 & x110 & x111 & x112))) | (x103 & (~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x101 | ~x102)));
  assign z75 = x004 & ~x006 & ((x101 & x102 & x103 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x104) | (x113 & x114 & x115 & x116 & x110 & x111 & x112 & x104 & x105 & x106 & x107 & x108 & x109))) | (x104 & (~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x101 | ~x102 | ~x103)));
  assign z76 = x004 & ((~x006 & ((x101 & x102 & x103 & x104 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x105) | (x105 & x106 & x107 & x108 & x109 & x110 & x111 & x112 & x113 & x114 & x115 & x116))) | (x105 & ((x005 & (~x103 | ~x104 | ~x101 | ~x102)) | ~x031 | ~x032 | x033 | ~x003 | ~x029 | ~x030)))) | (x003 & ~x005 & x029 & x030 & x031 & x032 & ~x033 & (~x105 | (x006 & (~x109 | ~x110 | ~x111 | ~x112 | ~x113 | ~x114 | ~x115 | ~x116 | ~x101 | ~x102 | ~x103 | ~x107 | ~x108 | ~x104 | ~x106)))));
  assign z77 = x004 & ~x006 & ((x105 & ((x109 & x110 & x111 & x112 & x113 & x114 & x115 & x116 & x101 & x102 & x103 & x107 & x108 & x104 & x106) | (x003 & x029 & x030 & x031 & x032 & ~x033 & ~x106 & (~x005 | (x103 & x104 & x101 & x102))))) | (x106 & ((x005 & (~x103 | ~x104 | ~x101 | ~x102)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x105)));
  assign z78 = x004 & ~x006 & ((x105 & x106 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x107 & (~x005 | (x103 & x104 & x101 & x102))) | (x113 & x114 & x115 & x116 & x110 & x111 & x112 & x101 & x102 & x103 & x108 & x109 & x104 & x107))) | (x107 & ((x005 & (~x103 | ~x104 | ~x101 | ~x102)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x105 | ~x106)));
  assign z79 = x004 & ~x006 & ((x105 & x106 & x107 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x108 & (~x005 | (x103 & x104 & x101 & x102))) | (x113 & x114 & x115 & x116 & x110 & x111 & x112 & x101 & x102 & x103 & x104 & x108 & x109))) | (x108 & ((x005 & (~x103 | ~x104 | ~x101 | ~x102)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x105 | ~x106 | ~x107)));
  assign z80 = x004 & ((((x003 & ~x005 & x006 & x029 & x032 & ~x033 & x030 & x031) | (x005 & ~x006 & x109)) & (~x105 | ~x106 | ~x107 | ~x108 | ~x103 | ~x104 | ~x101 | ~x102)) | (x003 & x029 & x030 & x031 & x032 & ~x033 & (~x005 | (x105 & x106 & x107 & x108 & x103 & x104 & x101 & x102)) & (~x109 | (x006 & (~x113 | ~x114 | ~x115 | ~x116 | ~x110 | ~x111 | ~x112)))) | (~x006 & x109 & (~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | (x101 & x102 & x103 & x104 & x105 & x106 & x107 & x113 & x114 & x115 & x116 & x111 & x112 & x108 & x110))));
  assign z81 = x004 & ~x006 & ((x109 & ((x101 & x102 & x103 & x104 & x105 & x106 & x107 & x113 & x114 & x115 & x116 & x111 & x112 & x108 & x110) | (x003 & x029 & x030 & x031 & x032 & ~x033 & ~x110 & (~x005 | (x105 & x106 & x107 & x108 & x103 & x104 & x101 & x102))))) | (x110 & ((x005 & (~x105 | ~x106 | ~x107 | ~x108 | ~x103 | ~x104 | ~x101 | ~x102)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x109)));
  assign z82 = x004 & ~x006 & ((x109 & x110 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x111 & (~x005 | (x105 & x106 & x107 & x108 & x103 & x104 & x101 & x102))) | (x101 & x102 & x103 & x104 & x105 & x106 & x107 & x113 & x114 & x115 & x116 & x108 & x111 & x112))) | (x111 & ((x005 & (~x105 | ~x106 | ~x107 | ~x108 | ~x103 | ~x104 | ~x101 | ~x102)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x109 | ~x110)));
  assign z83 = x004 & ~x006 & ((x109 & x110 & x111 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x112 & (~x005 | (x105 & x106 & x107 & x108 & x103 & x104 & x101 & x102))) | (x104 & x105 & x106 & x101 & x102 & x103 & x113 & x114 & x115 & x116 & x107 & x108 & x112))) | (x112 & ((x005 & (~x105 | ~x106 | ~x107 | ~x108 | ~x103 | ~x104 | ~x101 | ~x102)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x109 | ~x110 | ~x111)));
  assign z84 = x004 & ((~x006 & ((x101 & x102 & x103 & x104 & x105 & x106 & x107 & x108 & x109 & x110 & x111 & x112 & ((x113 & x114 & x115 & x116) | (x003 & x029 & x030 & x031 & x032 & ~x033 & ~x113))) | (x113 & (~x031 | ~x032 | x033 | ~x003 | ~x029 | ~x030 | (x005 & (~x104 | ~x105 | ~x106 | ~x101 | ~x102 | ~x103 | ~x110 | ~x111 | ~x112 | ~x107 | ~x108 | ~x109)))))) | (x003 & ~x005 & x029 & x030 & x031 & x032 & ~x033 & (~x113 | (x006 & (~x101 | ~x102 | ~x103 | ~x104 | ~x105 | ~x106 | ~x107 | ~x108 | ~x109 | ~x110 | ~x111 | ~x115 | ~x116 | ~x112 | ~x114)))));
  assign z85 = x004 & ~x006 & ((x113 & ((x101 & x102 & x103 & x104 & x105 & x106 & x107 & x108 & x109 & x110 & x111 & x115 & x116 & x112 & x114) | (x003 & x029 & x030 & x031 & x032 & ~x033 & ~x114 & (~x005 | (x104 & x105 & x106 & x101 & x102 & x103 & x110 & x111 & x112 & x107 & x108 & x109))))) | (x114 & ((x005 & (~x104 | ~x105 | ~x106 | ~x101 | ~x102 | ~x103 | ~x110 | ~x111 | ~x112 | ~x107 | ~x108 | ~x109)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x113)));
  assign z86 = x004 & ~x006 & ((x113 & x114 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x115 & (~x005 | (x104 & x105 & x106 & x101 & x102 & x103 & x110 & x111 & x112 & x107 & x108 & x109))) | (x101 & x102 & x103 & x104 & x105 & x106 & x107 & x108 & x109 & x110 & x111 & x112 & x115 & x116))) | (x115 & ((x005 & (~x104 | ~x105 | ~x106 | ~x101 | ~x102 | ~x103 | ~x110 | ~x111 | ~x112 | ~x107 | ~x108 | ~x109)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x113 | ~x114)));
  assign z87 = x004 & ~x006 & ((x113 & x114 & x115 & ((x003 & x029 & x030 & x031 & x032 & ~x033 & ~x116 & (~x005 | (x104 & x105 & x106 & x101 & x102 & x103 & x110 & x111 & x112 & x107 & x108 & x109))) | (x104 & x105 & x106 & x101 & x102 & x103 & x107 & x108 & x109 & x110 & x111 & x112 & x116))) | (x116 & ((x005 & (~x104 | ~x105 | ~x106 | ~x101 | ~x102 | ~x103 | ~x110 | ~x111 | ~x112 | ~x107 | ~x108 | ~x109)) | ~x003 | ~x029 | ~x030 | ~x031 | ~x032 | x033 | ~x113 | ~x114 | ~x115)));
  assign z29 = 1'b0;
  assign z30 = 1'b0;
  assign z31 = 1'b0;
endmodule